
module HighActiveRegionDetection_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module HighActiveRegionDetection_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module HighActiveRegionDetection_DW01_inc_2 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module HighActiveRegionDetection_DW01_inc_3 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module HighActiveRegionDetection_DW01_inc_4 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module HighActiveRegionDetection_DW01_inc_5 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module HighActiveRegionDetection_DW01_inc_6 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module HighActiveRegionDetection_DW01_inc_7 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module HighActiveRegionDetection_DW01_inc_8 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HADDX1 U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  HADDX1 U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1 U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(carry[24]), .SO(SUM[23]) );
  HADDX1 U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1 U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1 U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  INVX0 U1 ( .IN(A[0]), .QN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[31]), .IN2(A[31]), .Q(SUM[31]) );
endmodule


module HighActiveRegionDetection ( clk, In0, In1, In2, In3, In4, In5, In6, In7, 
        Trigger_out );
  input clk, In0, In1, In2, In3, In4, In5, In6, In7;
  output Trigger_out;
  wire   N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, N35, N36, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N75, N76, N77, N78, N79, N80, N81,
         N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95,
         N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N145, N146,
         N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157,
         N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168,
         N169, N170, N171, N172, N173, N174, N175, N176, N180, N181, N182,
         N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193,
         N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N215, N216, N217, N218,
         N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348,
         N349, N350, N351, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761;
  wire   [31:0] Clock_counter;
  wire   [31:0] In7_counter;
  wire   [31:0] In6_counter;
  wire   [31:0] In5_counter;
  wire   [31:0] In4_counter;
  wire   [31:0] In3_counter;
  wire   [31:0] In2_counter;
  wire   [31:0] In1_counter;
  wire   [31:0] In0_counter;

  HighActiveRegionDetection_DW01_inc_0 add_141 ( .A(Clock_counter), .SUM({N319, 
        N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, 
        N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, 
        N294, N293, N292, N291, N290, N289, N288}) );
  HighActiveRegionDetection_DW01_inc_1 add_129 ( .A(In0_counter), .SUM({N281, 
        N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, 
        N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, 
        N256, N255, N254, N253, N252, N251, N250}) );
  HighActiveRegionDetection_DW01_inc_2 add_120 ( .A(In1_counter), .SUM({N246, 
        N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, 
        N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, 
        N221, N220, N219, N218, N217, N216, N215}) );
  HighActiveRegionDetection_DW01_inc_3 add_111 ( .A(In2_counter), .SUM({N211, 
        N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, 
        N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, 
        N186, N185, N184, N183, N182, N181, N180}) );
  HighActiveRegionDetection_DW01_inc_4 add_102 ( .A(In3_counter), .SUM({N176, 
        N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, 
        N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, 
        N151, N150, N149, N148, N147, N146, N145}) );
  HighActiveRegionDetection_DW01_inc_5 add_93 ( .A(In4_counter), .SUM({N141, 
        N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, 
        N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, 
        N116, N115, N114, N113, N112, N111, N110}) );
  HighActiveRegionDetection_DW01_inc_6 add_84 ( .A(In5_counter), .SUM({N106, 
        N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, 
        N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, 
        N78, N77, N76, N75}) );
  HighActiveRegionDetection_DW01_inc_7 add_75 ( .A(In6_counter), .SUM({N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40}) );
  HighActiveRegionDetection_DW01_inc_8 add_66 ( .A(In7_counter), .SUM({N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, 
        N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, 
        N6, N5}) );
  DFFARX1 Clock_counter_reg_31_ ( .D(N351), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[31]), .QN(n759) );
  DFFARX1 In5_counter_reg_31_ ( .D(N106), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[31]), .QN(n610) );
  DFFARX1 In7_counter_reg_31_ ( .D(N36), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[31]), .QN(n594) );
  DFFARX1 In0_counter_reg_31_ ( .D(N281), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[31]), .QN(n578) );
  DFFARX1 In2_counter_reg_31_ ( .D(N211), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[31]), .QN(n562) );
  DFFARX1 In4_counter_reg_31_ ( .D(N141), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[31]), .QN(n546) );
  DFFARX1 In3_counter_reg_31_ ( .D(N176), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[31]), .QN(n545) );
  DFFARX1 In1_counter_reg_31_ ( .D(N246), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[31]), .QN(n529) );
  DFFARX1 In6_counter_reg_31_ ( .D(N71), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[31]), .QN(n513) );
  DFFARX1 Clock_counter_reg_1_ ( .D(N321), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[1]), .QN(n758) );
  DFFARX1 In5_counter_reg_2_ ( .D(N77), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[2]), .QN(n625) );
  DFFARX1 In5_counter_reg_3_ ( .D(N78), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[3]), .QN(n624) );
  DFFARX1 In5_counter_reg_8_ ( .D(N83), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[8]), .QN(n623) );
  DFFARX1 In5_counter_reg_9_ ( .D(N84), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[9]), .QN(n622) );
  DFFARX1 In5_counter_reg_10_ ( .D(N85), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[10]), .QN(n621) );
  DFFARX1 In5_counter_reg_14_ ( .D(N89), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[14]), .QN(n620) );
  DFFARX1 In5_counter_reg_15_ ( .D(N90), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[15]), .QN(n619) );
  DFFARX1 In5_counter_reg_16_ ( .D(N91), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[16]), .QN(n618) );
  DFFARX1 In5_counter_reg_17_ ( .D(N92), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[17]), .QN(n617) );
  DFFARX1 In5_counter_reg_21_ ( .D(N96), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[21]), .QN(n616) );
  DFFARX1 In5_counter_reg_22_ ( .D(N97), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[22]), .QN(n615) );
  DFFARX1 In5_counter_reg_23_ ( .D(N98), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[23]), .QN(n614) );
  DFFARX1 In5_counter_reg_27_ ( .D(N102), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[27]), .QN(n613) );
  DFFARX1 In5_counter_reg_28_ ( .D(N103), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[28]), .QN(n612) );
  DFFARX1 In5_counter_reg_29_ ( .D(N104), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[29]), .QN(n611) );
  DFFARX1 In7_counter_reg_2_ ( .D(N7), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[2]), .QN(n609) );
  DFFARX1 In7_counter_reg_3_ ( .D(N8), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[3]), .QN(n608) );
  DFFARX1 In7_counter_reg_8_ ( .D(N13), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[8]), .QN(n607) );
  DFFARX1 In7_counter_reg_9_ ( .D(N14), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[9]), .QN(n606) );
  DFFARX1 In7_counter_reg_10_ ( .D(N15), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[10]), .QN(n605) );
  DFFARX1 In7_counter_reg_14_ ( .D(N19), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[14]), .QN(n604) );
  DFFARX1 In7_counter_reg_15_ ( .D(N20), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[15]), .QN(n603) );
  DFFARX1 In7_counter_reg_16_ ( .D(N21), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[16]), .QN(n602) );
  DFFARX1 In7_counter_reg_17_ ( .D(N22), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[17]), .QN(n601) );
  DFFARX1 In7_counter_reg_21_ ( .D(N26), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[21]), .QN(n600) );
  DFFARX1 In7_counter_reg_22_ ( .D(N27), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[22]), .QN(n599) );
  DFFARX1 In7_counter_reg_23_ ( .D(N28), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[23]), .QN(n598) );
  DFFARX1 In7_counter_reg_27_ ( .D(N32), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[27]), .QN(n597) );
  DFFARX1 In7_counter_reg_28_ ( .D(N33), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[28]), .QN(n596) );
  DFFARX1 In7_counter_reg_29_ ( .D(N34), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[29]), .QN(n595) );
  DFFARX1 In0_counter_reg_2_ ( .D(N252), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[2]), .QN(n593) );
  DFFARX1 In0_counter_reg_3_ ( .D(N253), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[3]), .QN(n592) );
  DFFARX1 In0_counter_reg_8_ ( .D(N258), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[8]), .QN(n591) );
  DFFARX1 In0_counter_reg_9_ ( .D(N259), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[9]), .QN(n590) );
  DFFARX1 In0_counter_reg_10_ ( .D(N260), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[10]), .QN(n589) );
  DFFARX1 In0_counter_reg_14_ ( .D(N264), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[14]), .QN(n588) );
  DFFARX1 In0_counter_reg_15_ ( .D(N265), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[15]), .QN(n587) );
  DFFARX1 In0_counter_reg_16_ ( .D(N266), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[16]), .QN(n586) );
  DFFARX1 In0_counter_reg_17_ ( .D(N267), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[17]), .QN(n585) );
  DFFARX1 In0_counter_reg_21_ ( .D(N271), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[21]), .QN(n584) );
  DFFARX1 In0_counter_reg_22_ ( .D(N272), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[22]), .QN(n583) );
  DFFARX1 In0_counter_reg_23_ ( .D(N273), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[23]), .QN(n582) );
  DFFARX1 In0_counter_reg_27_ ( .D(N277), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[27]), .QN(n581) );
  DFFARX1 In0_counter_reg_28_ ( .D(N278), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[28]), .QN(n580) );
  DFFARX1 In0_counter_reg_29_ ( .D(N279), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[29]), .QN(n579) );
  DFFARX1 In2_counter_reg_2_ ( .D(N182), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[2]), .QN(n577) );
  DFFARX1 In2_counter_reg_3_ ( .D(N183), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[3]), .QN(n576) );
  DFFARX1 In2_counter_reg_8_ ( .D(N188), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[8]), .QN(n575) );
  DFFARX1 In2_counter_reg_9_ ( .D(N189), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[9]), .QN(n574) );
  DFFARX1 In2_counter_reg_10_ ( .D(N190), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[10]), .QN(n573) );
  DFFARX1 In2_counter_reg_14_ ( .D(N194), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[14]), .QN(n572) );
  DFFARX1 In2_counter_reg_15_ ( .D(N195), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[15]), .QN(n571) );
  DFFARX1 In2_counter_reg_16_ ( .D(N196), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[16]), .QN(n570) );
  DFFARX1 In2_counter_reg_17_ ( .D(N197), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[17]), .QN(n569) );
  DFFARX1 In2_counter_reg_21_ ( .D(N201), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[21]), .QN(n568) );
  DFFARX1 In2_counter_reg_22_ ( .D(N202), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[22]), .QN(n567) );
  DFFARX1 In2_counter_reg_23_ ( .D(N203), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[23]), .QN(n566) );
  DFFARX1 In2_counter_reg_27_ ( .D(N207), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[27]), .QN(n565) );
  DFFARX1 In2_counter_reg_28_ ( .D(N208), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[28]), .QN(n564) );
  DFFARX1 In2_counter_reg_29_ ( .D(N209), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[29]), .QN(n563) );
  DFFARX1 In4_counter_reg_2_ ( .D(N112), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[2]), .QN(n561) );
  DFFARX1 In4_counter_reg_3_ ( .D(N113), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[3]), .QN(n560) );
  DFFARX1 In4_counter_reg_8_ ( .D(N118), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[8]), .QN(n559) );
  DFFARX1 In4_counter_reg_9_ ( .D(N119), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[9]), .QN(n558) );
  DFFARX1 In4_counter_reg_10_ ( .D(N120), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[10]), .QN(n557) );
  DFFARX1 In4_counter_reg_14_ ( .D(N124), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[14]), .QN(n556) );
  DFFARX1 In4_counter_reg_15_ ( .D(N125), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[15]), .QN(n555) );
  DFFARX1 In4_counter_reg_16_ ( .D(N126), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[16]), .QN(n554) );
  DFFARX1 In4_counter_reg_17_ ( .D(N127), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[17]), .QN(n553) );
  DFFARX1 In4_counter_reg_21_ ( .D(N131), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[21]), .QN(n552) );
  DFFARX1 In4_counter_reg_22_ ( .D(N132), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[22]), .QN(n551) );
  DFFARX1 In4_counter_reg_23_ ( .D(N133), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[23]), .QN(n550) );
  DFFARX1 In4_counter_reg_27_ ( .D(N137), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[27]), .QN(n549) );
  DFFARX1 In4_counter_reg_28_ ( .D(N138), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[28]), .QN(n548) );
  DFFARX1 In4_counter_reg_29_ ( .D(N139), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[29]), .QN(n547) );
  DFFARX1 In3_counter_reg_2_ ( .D(N147), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[2]), .QN(n544) );
  DFFARX1 In3_counter_reg_3_ ( .D(N148), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[3]), .QN(n543) );
  DFFARX1 In3_counter_reg_9_ ( .D(N154), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[9]), .QN(n542) );
  DFFARX1 In3_counter_reg_10_ ( .D(N155), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[10]), .QN(n541) );
  DFFARX1 In3_counter_reg_11_ ( .D(N156), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[11]), .QN(n540) );
  DFFARX1 In3_counter_reg_15_ ( .D(N160), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[15]), .QN(n539) );
  DFFARX1 In3_counter_reg_16_ ( .D(N161), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[16]), .QN(n538) );
  DFFARX1 In3_counter_reg_17_ ( .D(N162), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[17]), .QN(n537) );
  DFFARX1 In3_counter_reg_18_ ( .D(N163), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[18]), .QN(n536) );
  DFFARX1 In3_counter_reg_22_ ( .D(N167), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[22]), .QN(n535) );
  DFFARX1 In3_counter_reg_23_ ( .D(N168), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[23]), .QN(n534) );
  DFFARX1 In3_counter_reg_24_ ( .D(N169), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[24]), .QN(n533) );
  DFFARX1 In3_counter_reg_28_ ( .D(N173), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[28]), .QN(n532) );
  DFFARX1 In3_counter_reg_29_ ( .D(N174), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[29]), .QN(n531) );
  DFFARX1 In3_counter_reg_30_ ( .D(N175), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[30]), .QN(n530) );
  DFFARX1 In1_counter_reg_2_ ( .D(N217), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[2]), .QN(n528) );
  DFFARX1 In1_counter_reg_3_ ( .D(N218), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[3]), .QN(n527) );
  DFFARX1 In1_counter_reg_9_ ( .D(N224), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[9]), .QN(n526) );
  DFFARX1 In1_counter_reg_10_ ( .D(N225), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[10]), .QN(n525) );
  DFFARX1 In1_counter_reg_11_ ( .D(N226), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[11]), .QN(n524) );
  DFFARX1 In1_counter_reg_15_ ( .D(N230), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[15]), .QN(n523) );
  DFFARX1 In1_counter_reg_16_ ( .D(N231), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[16]), .QN(n522) );
  DFFARX1 In1_counter_reg_17_ ( .D(N232), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[17]), .QN(n521) );
  DFFARX1 In1_counter_reg_18_ ( .D(N233), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[18]), .QN(n520) );
  DFFARX1 In1_counter_reg_22_ ( .D(N237), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[22]), .QN(n519) );
  DFFARX1 In1_counter_reg_23_ ( .D(N238), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[23]), .QN(n518) );
  DFFARX1 In1_counter_reg_24_ ( .D(N239), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[24]), .QN(n517) );
  DFFARX1 In1_counter_reg_28_ ( .D(N243), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[28]), .QN(n516) );
  DFFARX1 In1_counter_reg_29_ ( .D(N244), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[29]), .QN(n515) );
  DFFARX1 In1_counter_reg_30_ ( .D(N245), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[30]), .QN(n514) );
  DFFARX1 Clock_counter_reg_27_ ( .D(N347), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[27]), .QN(n757) );
  DFFARX1 Clock_counter_reg_26_ ( .D(N346), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[26]), .QN(n756) );
  DFFARX1 Clock_counter_reg_25_ ( .D(N345), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[25]), .QN(n755) );
  DFFARX1 Clock_counter_reg_21_ ( .D(N341), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[21]), .QN(n754) );
  DFFARX1 Clock_counter_reg_20_ ( .D(N340), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[20]), .QN(n753) );
  DFFARX1 Clock_counter_reg_19_ ( .D(N339), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[19]), .QN(n752) );
  DFFARX1 Clock_counter_reg_15_ ( .D(N335), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[15]), .QN(n751) );
  DFFARX1 Clock_counter_reg_14_ ( .D(N334), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[14]), .QN(n750) );
  DFFARX1 Clock_counter_reg_13_ ( .D(N333), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[13]), .QN(n749) );
  DFFARX1 Clock_counter_reg_9_ ( .D(N329), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[9]), .QN(n748) );
  DFFARX1 Clock_counter_reg_8_ ( .D(N328), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[8]), .QN(n747) );
  DFFARX1 Clock_counter_reg_7_ ( .D(N327), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[7]), .QN(n746) );
  DFFARX1 Clock_counter_reg_3_ ( .D(N323), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[3]), .QN() );
  DFFARX1 Clock_counter_reg_2_ ( .D(N322), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[2]), .QN() );
  DFFARX1 In6_counter_reg_2_ ( .D(N42), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[2]), .QN(n512) );
  DFFARX1 In6_counter_reg_3_ ( .D(N43), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[3]), .QN(n511) );
  DFFARX1 In6_counter_reg_9_ ( .D(N49), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[9]), .QN(n510) );
  DFFARX1 In6_counter_reg_10_ ( .D(N50), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[10]), .QN(n509) );
  DFFARX1 In6_counter_reg_11_ ( .D(N51), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[11]), .QN(n508) );
  DFFARX1 In6_counter_reg_15_ ( .D(N55), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[15]), .QN(n507) );
  DFFARX1 In6_counter_reg_16_ ( .D(N56), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[16]), .QN(n506) );
  DFFARX1 In6_counter_reg_17_ ( .D(N57), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[17]), .QN(n505) );
  DFFARX1 In6_counter_reg_18_ ( .D(N58), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[18]), .QN(n504) );
  DFFARX1 In6_counter_reg_22_ ( .D(N62), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[22]), .QN(n503) );
  DFFARX1 In6_counter_reg_23_ ( .D(N63), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[23]), .QN(n502) );
  DFFARX1 In6_counter_reg_24_ ( .D(N64), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[24]), .QN(n501) );
  DFFARX1 In6_counter_reg_28_ ( .D(N68), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[28]), .QN(n500) );
  DFFARX1 In6_counter_reg_29_ ( .D(N69), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[29]), .QN(n499) );
  DFFARX1 In6_counter_reg_30_ ( .D(N70), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[30]), .QN(n498) );
  DFFARX1 Clock_counter_reg_4_ ( .D(N324), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[4]), .QN() );
  DFFARX1 In5_counter_reg_1_ ( .D(N76), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[1]), .QN() );
  DFFARX1 In7_counter_reg_1_ ( .D(N6), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[1]), .QN() );
  DFFARX1 In0_counter_reg_1_ ( .D(N251), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[1]), .QN() );
  DFFARX1 In2_counter_reg_1_ ( .D(N181), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[1]), .QN() );
  DFFARX1 In4_counter_reg_1_ ( .D(N111), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[1]), .QN() );
  DFFARX1 In3_counter_reg_1_ ( .D(N146), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[1]), .QN() );
  DFFARX1 In1_counter_reg_1_ ( .D(N216), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[1]), .QN() );
  DFFARX1 In6_counter_reg_1_ ( .D(N41), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[1]), .QN() );
  DFFARX1 Clock_counter_reg_5_ ( .D(N325), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[5]), .QN() );
  DFFARX1 Clock_counter_reg_6_ ( .D(N326), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[6]), .QN() );
  DFFARX1 In5_counter_reg_5_ ( .D(N80), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[5]), .QN() );
  DFFARX1 In7_counter_reg_5_ ( .D(N10), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[5]), .QN() );
  DFFARX1 In0_counter_reg_5_ ( .D(N255), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[5]), .QN() );
  DFFARX1 In2_counter_reg_5_ ( .D(N185), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[5]), .QN() );
  DFFARX1 In4_counter_reg_5_ ( .D(N115), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[5]), .QN() );
  DFFARX1 In3_counter_reg_5_ ( .D(N150), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[5]), .QN() );
  DFFARX1 In1_counter_reg_5_ ( .D(N220), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[5]), .QN() );
  DFFARX1 In6_counter_reg_5_ ( .D(N45), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[5]), .QN() );
  DFFARX1 In5_counter_reg_4_ ( .D(N79), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[4]), .QN() );
  DFFARX1 In7_counter_reg_4_ ( .D(N9), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[4]), .QN() );
  DFFARX1 In0_counter_reg_4_ ( .D(N254), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[4]), .QN() );
  DFFARX1 In2_counter_reg_4_ ( .D(N184), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[4]), .QN() );
  DFFARX1 In4_counter_reg_4_ ( .D(N114), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[4]), .QN() );
  DFFARX1 In3_counter_reg_4_ ( .D(N149), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[4]), .QN() );
  DFFARX1 In1_counter_reg_4_ ( .D(N219), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[4]), .QN() );
  DFFARX1 In6_counter_reg_4_ ( .D(N44), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[4]), .QN() );
  DFFARX1 In5_counter_reg_30_ ( .D(N105), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[30]), .QN() );
  DFFARX1 In5_counter_reg_11_ ( .D(N86), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[11]), .QN() );
  DFFARX1 In5_counter_reg_18_ ( .D(N93), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[18]), .QN() );
  DFFARX1 In5_counter_reg_24_ ( .D(N99), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[24]), .QN() );
  DFFARX1 In7_counter_reg_30_ ( .D(N35), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[30]), .QN() );
  DFFARX1 In7_counter_reg_11_ ( .D(N16), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[11]), .QN() );
  DFFARX1 In7_counter_reg_18_ ( .D(N23), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[18]), .QN() );
  DFFARX1 In7_counter_reg_24_ ( .D(N29), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[24]), .QN() );
  DFFARX1 In0_counter_reg_30_ ( .D(N280), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[30]), .QN() );
  DFFARX1 In0_counter_reg_11_ ( .D(N261), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[11]), .QN() );
  DFFARX1 In0_counter_reg_18_ ( .D(N268), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[18]), .QN() );
  DFFARX1 In0_counter_reg_24_ ( .D(N274), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[24]), .QN() );
  DFFARX1 In2_counter_reg_30_ ( .D(N210), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[30]), .QN() );
  DFFARX1 In2_counter_reg_11_ ( .D(N191), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[11]), .QN() );
  DFFARX1 In2_counter_reg_18_ ( .D(N198), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[18]), .QN() );
  DFFARX1 In2_counter_reg_24_ ( .D(N204), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[24]), .QN() );
  DFFARX1 In4_counter_reg_30_ ( .D(N140), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[30]), .QN() );
  DFFARX1 In4_counter_reg_11_ ( .D(N121), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[11]), .QN() );
  DFFARX1 In4_counter_reg_18_ ( .D(N128), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[18]), .QN() );
  DFFARX1 In4_counter_reg_24_ ( .D(N134), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[24]), .QN() );
  DFFARX1 In3_counter_reg_6_ ( .D(N151), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[6]), .QN() );
  DFFARX1 In3_counter_reg_12_ ( .D(N157), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[12]), .QN() );
  DFFARX1 In3_counter_reg_19_ ( .D(N164), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[19]), .QN() );
  DFFARX1 In3_counter_reg_25_ ( .D(N170), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[25]), .QN() );
  DFFARX1 In1_counter_reg_6_ ( .D(N221), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[6]), .QN() );
  DFFARX1 In1_counter_reg_12_ ( .D(N227), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[12]), .QN() );
  DFFARX1 In1_counter_reg_19_ ( .D(N234), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[19]), .QN() );
  DFFARX1 In1_counter_reg_25_ ( .D(N240), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[25]), .QN() );
  DFFARX1 Clock_counter_reg_30_ ( .D(N350), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[30]), .QN() );
  DFFARX1 Clock_counter_reg_24_ ( .D(N344), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[24]), .QN() );
  DFFARX1 Clock_counter_reg_18_ ( .D(N338), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[18]), .QN() );
  DFFARX1 Clock_counter_reg_12_ ( .D(N332), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[12]), .QN() );
  DFFARX1 In6_counter_reg_6_ ( .D(N46), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[6]), .QN() );
  DFFARX1 In6_counter_reg_12_ ( .D(N52), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[12]), .QN() );
  DFFARX1 In6_counter_reg_19_ ( .D(N59), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[19]), .QN() );
  DFFARX1 In6_counter_reg_25_ ( .D(N65), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[25]), .QN() );
  DFFARX1 In5_counter_reg_7_ ( .D(N82), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[7]), .QN() );
  DFFARX1 In5_counter_reg_13_ ( .D(N88), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[13]), .QN() );
  DFFARX1 In5_counter_reg_20_ ( .D(N95), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[20]), .QN() );
  DFFARX1 In5_counter_reg_26_ ( .D(N101), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[26]), .QN() );
  DFFARX1 In7_counter_reg_7_ ( .D(N12), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[7]), .QN() );
  DFFARX1 In7_counter_reg_13_ ( .D(N18), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[13]), .QN() );
  DFFARX1 In7_counter_reg_20_ ( .D(N25), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[20]), .QN() );
  DFFARX1 In7_counter_reg_26_ ( .D(N31), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[26]), .QN() );
  DFFARX1 In0_counter_reg_7_ ( .D(N257), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[7]), .QN() );
  DFFARX1 In0_counter_reg_13_ ( .D(N263), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[13]), .QN() );
  DFFARX1 In0_counter_reg_20_ ( .D(N270), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[20]), .QN() );
  DFFARX1 In0_counter_reg_26_ ( .D(N276), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[26]), .QN() );
  DFFARX1 In2_counter_reg_7_ ( .D(N187), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[7]), .QN() );
  DFFARX1 In2_counter_reg_13_ ( .D(N193), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[13]), .QN() );
  DFFARX1 In2_counter_reg_20_ ( .D(N200), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[20]), .QN() );
  DFFARX1 In2_counter_reg_26_ ( .D(N206), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[26]), .QN() );
  DFFARX1 In4_counter_reg_7_ ( .D(N117), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[7]), .QN() );
  DFFARX1 In4_counter_reg_13_ ( .D(N123), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[13]), .QN() );
  DFFARX1 In4_counter_reg_20_ ( .D(N130), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[20]), .QN() );
  DFFARX1 In4_counter_reg_26_ ( .D(N136), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[26]), .QN() );
  DFFARX1 In3_counter_reg_8_ ( .D(N153), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[8]), .QN() );
  DFFARX1 In3_counter_reg_14_ ( .D(N159), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[14]), .QN() );
  DFFARX1 In3_counter_reg_21_ ( .D(N166), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[21]), .QN() );
  DFFARX1 In3_counter_reg_27_ ( .D(N172), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[27]), .QN() );
  DFFARX1 In1_counter_reg_8_ ( .D(N223), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[8]), .QN() );
  DFFARX1 In1_counter_reg_14_ ( .D(N229), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[14]), .QN() );
  DFFARX1 In1_counter_reg_21_ ( .D(N236), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[21]), .QN() );
  DFFARX1 In1_counter_reg_27_ ( .D(N242), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[27]), .QN() );
  DFFARX1 Clock_counter_reg_28_ ( .D(N348), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[28]), .QN() );
  DFFARX1 Clock_counter_reg_22_ ( .D(N342), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[22]), .QN() );
  DFFARX1 Clock_counter_reg_16_ ( .D(N336), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[16]), .QN() );
  DFFARX1 Clock_counter_reg_10_ ( .D(N330), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[10]), .QN() );
  DFFARX1 In6_counter_reg_8_ ( .D(N48), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[8]), .QN() );
  DFFARX1 In6_counter_reg_14_ ( .D(N54), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[14]), .QN() );
  DFFARX1 In6_counter_reg_21_ ( .D(N61), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[21]), .QN() );
  DFFARX1 In6_counter_reg_27_ ( .D(N67), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[27]), .QN() );
  DFFARX1 In5_counter_reg_6_ ( .D(N81), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[6]), .QN() );
  DFFARX1 In5_counter_reg_12_ ( .D(N87), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[12]), .QN() );
  DFFARX1 In5_counter_reg_19_ ( .D(N94), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[19]), .QN() );
  DFFARX1 In5_counter_reg_25_ ( .D(N100), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[25]), .QN() );
  DFFARX1 In7_counter_reg_6_ ( .D(N11), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[6]), .QN() );
  DFFARX1 In7_counter_reg_12_ ( .D(N17), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[12]), .QN() );
  DFFARX1 In7_counter_reg_19_ ( .D(N24), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[19]), .QN() );
  DFFARX1 In7_counter_reg_25_ ( .D(N30), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[25]), .QN() );
  DFFARX1 In0_counter_reg_6_ ( .D(N256), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[6]), .QN() );
  DFFARX1 In0_counter_reg_12_ ( .D(N262), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[12]), .QN() );
  DFFARX1 In0_counter_reg_19_ ( .D(N269), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[19]), .QN() );
  DFFARX1 In0_counter_reg_25_ ( .D(N275), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[25]), .QN() );
  DFFARX1 In2_counter_reg_6_ ( .D(N186), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[6]), .QN() );
  DFFARX1 In2_counter_reg_12_ ( .D(N192), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[12]), .QN() );
  DFFARX1 In2_counter_reg_19_ ( .D(N199), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[19]), .QN() );
  DFFARX1 In2_counter_reg_25_ ( .D(N205), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[25]), .QN() );
  DFFARX1 In4_counter_reg_6_ ( .D(N116), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[6]), .QN() );
  DFFARX1 In4_counter_reg_12_ ( .D(N122), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[12]), .QN() );
  DFFARX1 In4_counter_reg_19_ ( .D(N129), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[19]), .QN() );
  DFFARX1 In4_counter_reg_25_ ( .D(N135), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[25]), .QN() );
  DFFARX1 In3_counter_reg_7_ ( .D(N152), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[7]), .QN() );
  DFFARX1 In3_counter_reg_13_ ( .D(N158), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[13]), .QN() );
  DFFARX1 In3_counter_reg_20_ ( .D(N165), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[20]), .QN() );
  DFFARX1 In3_counter_reg_26_ ( .D(N171), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[26]), .QN() );
  DFFARX1 In1_counter_reg_7_ ( .D(N222), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[7]), .QN() );
  DFFARX1 In1_counter_reg_13_ ( .D(N228), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[13]), .QN() );
  DFFARX1 In1_counter_reg_20_ ( .D(N235), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[20]), .QN() );
  DFFARX1 In1_counter_reg_26_ ( .D(N241), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[26]), .QN() );
  DFFARX1 Clock_counter_reg_29_ ( .D(N349), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[29]), .QN() );
  DFFARX1 Clock_counter_reg_23_ ( .D(N343), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[23]), .QN() );
  DFFARX1 Clock_counter_reg_17_ ( .D(N337), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[17]), .QN() );
  DFFARX1 Clock_counter_reg_11_ ( .D(N331), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[11]), .QN() );
  DFFARX1 In6_counter_reg_7_ ( .D(N47), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[7]), .QN() );
  DFFARX1 In6_counter_reg_13_ ( .D(N53), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[13]), .QN() );
  DFFARX1 In6_counter_reg_20_ ( .D(N60), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[20]), .QN() );
  DFFARX1 In6_counter_reg_26_ ( .D(N66), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[26]), .QN() );
  DFFARX1 Clock_counter_reg_0_ ( .D(N320), .CLK(clk), .RSTB(n761), .Q(
        Clock_counter[0]), .QN(n760) );
  DFFARX1 In5_counter_reg_0_ ( .D(N75), .CLK(In5), .RSTB(n761), .Q(
        In5_counter[0]), .QN() );
  DFFARX1 In7_counter_reg_0_ ( .D(N5), .CLK(In7), .RSTB(n761), .Q(
        In7_counter[0]), .QN() );
  DFFARX1 In0_counter_reg_0_ ( .D(N250), .CLK(In0), .RSTB(n761), .Q(
        In0_counter[0]), .QN() );
  DFFARX1 In2_counter_reg_0_ ( .D(N180), .CLK(In2), .RSTB(n761), .Q(
        In2_counter[0]), .QN() );
  DFFARX1 In4_counter_reg_0_ ( .D(N110), .CLK(In4), .RSTB(n761), .Q(
        In4_counter[0]), .QN() );
  DFFARX1 In3_counter_reg_0_ ( .D(N145), .CLK(In3), .RSTB(n761), .Q(
        In3_counter[0]), .QN() );
  DFFARX1 In1_counter_reg_0_ ( .D(N215), .CLK(In1), .RSTB(n761), .Q(
        In1_counter[0]), .QN() );
  DFFARX1 In6_counter_reg_0_ ( .D(N40), .CLK(In6), .RSTB(n761), .Q(
        In6_counter[0]), .QN() );
  OA21X1 U64 ( .IN1(n626), .IN2(n627), .IN3(n628), .Q(n761) );
  INVX0 U65 ( .IN(n629), .QN(n628) );
  OR4X1 U66 ( .IN1(In1), .IN2(In0), .IN3(In3), .IN4(In2), .Q(n627) );
  OR4X1 U67 ( .IN1(In5), .IN2(In4), .IN3(In7), .IN4(In6), .Q(n626) );
  NOR4X0 U68 ( .IN1(n630), .IN2(n631), .IN3(n632), .IN4(n633), .QN(Trigger_out) );
  NAND4X0 U69 ( .IN1(n610), .IN2(n594), .IN3(n578), .IN4(n562), .QN(n633) );
  NAND4X0 U70 ( .IN1(n546), .IN2(n545), .IN3(n529), .IN4(n513), .QN(n632) );
  NAND4X0 U71 ( .IN1(n634), .IN2(n635), .IN3(n636), .IN4(n637), .QN(n631) );
  NAND4X0 U72 ( .IN1(n638), .IN2(n639), .IN3(n640), .IN4(n641), .QN(n637) );
  NOR4X0 U73 ( .IN1(n642), .IN2(In0_counter[24]), .IN3(In0_counter[26]), .IN4(
        In0_counter[25]), .QN(n641) );
  NAND4X0 U74 ( .IN1(n581), .IN2(n580), .IN3(n579), .IN4(n643), .QN(n642) );
  NAND3X0 U75 ( .IN1(In0_counter[5]), .IN2(In0_counter[4]), .IN3(n644), .QN(
        n643) );
  NAND3X0 U76 ( .IN1(n592), .IN2(n645), .IN3(n593), .QN(n644) );
  NAND2X0 U77 ( .IN1(In0_counter[1]), .IN2(In0_counter[0]), .QN(n645) );
  NOR4X0 U78 ( .IN1(n646), .IN2(In0_counter[18]), .IN3(In0_counter[20]), .IN4(
        In0_counter[19]), .QN(n640) );
  NAND3X0 U79 ( .IN1(n583), .IN2(n582), .IN3(n584), .QN(n646) );
  NOR4X0 U80 ( .IN1(n647), .IN2(In0_counter[11]), .IN3(In0_counter[13]), .IN4(
        In0_counter[12]), .QN(n639) );
  NAND4X0 U81 ( .IN1(n588), .IN2(n587), .IN3(n586), .IN4(n585), .QN(n647) );
  NOR4X0 U82 ( .IN1(n648), .IN2(In0_counter[30]), .IN3(In0_counter[7]), .IN4(
        In0_counter[6]), .QN(n638) );
  NAND3X0 U83 ( .IN1(n590), .IN2(n589), .IN3(n591), .QN(n648) );
  NAND4X0 U84 ( .IN1(n649), .IN2(n650), .IN3(n651), .IN4(n652), .QN(n636) );
  NOR4X0 U85 ( .IN1(n653), .IN2(In2_counter[24]), .IN3(In2_counter[26]), .IN4(
        In2_counter[25]), .QN(n652) );
  NAND4X0 U86 ( .IN1(n565), .IN2(n564), .IN3(n563), .IN4(n654), .QN(n653) );
  NAND3X0 U87 ( .IN1(In2_counter[5]), .IN2(In2_counter[4]), .IN3(n655), .QN(
        n654) );
  NAND3X0 U88 ( .IN1(n576), .IN2(n656), .IN3(n577), .QN(n655) );
  NAND2X0 U89 ( .IN1(In2_counter[1]), .IN2(In2_counter[0]), .QN(n656) );
  NOR4X0 U90 ( .IN1(n657), .IN2(In2_counter[18]), .IN3(In2_counter[20]), .IN4(
        In2_counter[19]), .QN(n651) );
  NAND3X0 U91 ( .IN1(n567), .IN2(n566), .IN3(n568), .QN(n657) );
  NOR4X0 U92 ( .IN1(n658), .IN2(In2_counter[11]), .IN3(In2_counter[13]), .IN4(
        In2_counter[12]), .QN(n650) );
  NAND4X0 U93 ( .IN1(n572), .IN2(n571), .IN3(n570), .IN4(n569), .QN(n658) );
  NOR4X0 U94 ( .IN1(n659), .IN2(In2_counter[30]), .IN3(In2_counter[7]), .IN4(
        In2_counter[6]), .QN(n649) );
  NAND3X0 U95 ( .IN1(n574), .IN2(n573), .IN3(n575), .QN(n659) );
  NAND4X0 U96 ( .IN1(n660), .IN2(n661), .IN3(n662), .IN4(n663), .QN(n635) );
  NOR4X0 U97 ( .IN1(n664), .IN2(In3_counter[25]), .IN3(In3_counter[27]), .IN4(
        In3_counter[26]), .QN(n663) );
  NAND4X0 U98 ( .IN1(n532), .IN2(n531), .IN3(n530), .IN4(n665), .QN(n664) );
  NAND3X0 U99 ( .IN1(In3_counter[5]), .IN2(In3_counter[4]), .IN3(n666), .QN(
        n665) );
  NAND3X0 U100 ( .IN1(n543), .IN2(n667), .IN3(n544), .QN(n666) );
  NAND2X0 U101 ( .IN1(In3_counter[1]), .IN2(In3_counter[0]), .QN(n667) );
  NOR4X0 U102 ( .IN1(n668), .IN2(In3_counter[19]), .IN3(In3_counter[21]), 
        .IN4(In3_counter[20]), .QN(n662) );
  NAND3X0 U103 ( .IN1(n534), .IN2(n533), .IN3(n535), .QN(n668) );
  NOR4X0 U104 ( .IN1(n669), .IN2(In3_counter[12]), .IN3(In3_counter[14]), 
        .IN4(In3_counter[13]), .QN(n661) );
  NAND4X0 U105 ( .IN1(n539), .IN2(n538), .IN3(n537), .IN4(n536), .QN(n669) );
  NOR4X0 U106 ( .IN1(n670), .IN2(In3_counter[6]), .IN3(In3_counter[8]), .IN4(
        In3_counter[7]), .QN(n660) );
  NAND3X0 U107 ( .IN1(n541), .IN2(n540), .IN3(n542), .QN(n670) );
  OAI21X1 U108 ( .IN1(n671), .IN2(n672), .IN3(n759), .QN(n634) );
  OA21X1 U109 ( .IN1(Clock_counter[2]), .IN2(Clock_counter[3]), .IN3(n673), 
        .Q(n671) );
  NAND3X0 U110 ( .IN1(n674), .IN2(n675), .IN3(n676), .QN(n630) );
  AND3X1 U111 ( .IN1(n677), .IN2(n678), .IN3(n679), .Q(n676) );
  NAND4X0 U112 ( .IN1(n680), .IN2(n681), .IN3(n682), .IN4(n683), .QN(n679) );
  NOR4X0 U113 ( .IN1(n684), .IN2(In5_counter[24]), .IN3(In5_counter[26]), 
        .IN4(In5_counter[25]), .QN(n683) );
  NAND4X0 U114 ( .IN1(n613), .IN2(n612), .IN3(n611), .IN4(n685), .QN(n684) );
  NAND3X0 U115 ( .IN1(In5_counter[5]), .IN2(In5_counter[4]), .IN3(n686), .QN(
        n685) );
  NAND3X0 U116 ( .IN1(n624), .IN2(n687), .IN3(n625), .QN(n686) );
  NAND2X0 U117 ( .IN1(In5_counter[1]), .IN2(In5_counter[0]), .QN(n687) );
  NOR4X0 U118 ( .IN1(n688), .IN2(In5_counter[18]), .IN3(In5_counter[20]), 
        .IN4(In5_counter[19]), .QN(n682) );
  NAND3X0 U119 ( .IN1(n615), .IN2(n614), .IN3(n616), .QN(n688) );
  NOR4X0 U120 ( .IN1(n689), .IN2(In5_counter[11]), .IN3(In5_counter[13]), 
        .IN4(In5_counter[12]), .QN(n681) );
  NAND4X0 U121 ( .IN1(n620), .IN2(n619), .IN3(n618), .IN4(n617), .QN(n689) );
  NOR4X0 U122 ( .IN1(n690), .IN2(In5_counter[30]), .IN3(In5_counter[7]), .IN4(
        In5_counter[6]), .QN(n680) );
  NAND3X0 U123 ( .IN1(n622), .IN2(n621), .IN3(n623), .QN(n690) );
  NAND4X0 U124 ( .IN1(n691), .IN2(n692), .IN3(n693), .IN4(n694), .QN(n678) );
  NOR4X0 U125 ( .IN1(n695), .IN2(In7_counter[24]), .IN3(In7_counter[26]), 
        .IN4(In7_counter[25]), .QN(n694) );
  NAND4X0 U126 ( .IN1(n597), .IN2(n596), .IN3(n595), .IN4(n696), .QN(n695) );
  NAND3X0 U127 ( .IN1(In7_counter[5]), .IN2(In7_counter[4]), .IN3(n697), .QN(
        n696) );
  NAND3X0 U128 ( .IN1(n608), .IN2(n698), .IN3(n609), .QN(n697) );
  NAND2X0 U129 ( .IN1(In7_counter[1]), .IN2(In7_counter[0]), .QN(n698) );
  NOR4X0 U130 ( .IN1(n699), .IN2(In7_counter[18]), .IN3(In7_counter[20]), 
        .IN4(In7_counter[19]), .QN(n693) );
  NAND3X0 U131 ( .IN1(n599), .IN2(n598), .IN3(n600), .QN(n699) );
  NOR4X0 U132 ( .IN1(n700), .IN2(In7_counter[11]), .IN3(In7_counter[13]), 
        .IN4(In7_counter[12]), .QN(n692) );
  NAND4X0 U133 ( .IN1(n604), .IN2(n603), .IN3(n602), .IN4(n601), .QN(n700) );
  NOR4X0 U134 ( .IN1(n701), .IN2(In7_counter[30]), .IN3(In7_counter[7]), .IN4(
        In7_counter[6]), .QN(n691) );
  NAND3X0 U135 ( .IN1(n606), .IN2(n605), .IN3(n607), .QN(n701) );
  NAND4X0 U136 ( .IN1(n702), .IN2(n703), .IN3(n704), .IN4(n705), .QN(n677) );
  NOR4X0 U137 ( .IN1(n706), .IN2(In6_counter[25]), .IN3(In6_counter[27]), 
        .IN4(In6_counter[26]), .QN(n705) );
  NAND4X0 U138 ( .IN1(n500), .IN2(n499), .IN3(n498), .IN4(n707), .QN(n706) );
  NAND3X0 U139 ( .IN1(In6_counter[5]), .IN2(In6_counter[4]), .IN3(n708), .QN(
        n707) );
  NAND3X0 U140 ( .IN1(n511), .IN2(n709), .IN3(n512), .QN(n708) );
  NAND2X0 U141 ( .IN1(In6_counter[1]), .IN2(In6_counter[0]), .QN(n709) );
  NOR4X0 U142 ( .IN1(n710), .IN2(In6_counter[19]), .IN3(In6_counter[21]), 
        .IN4(In6_counter[20]), .QN(n704) );
  NAND3X0 U143 ( .IN1(n502), .IN2(n501), .IN3(n503), .QN(n710) );
  NOR4X0 U144 ( .IN1(n711), .IN2(In6_counter[12]), .IN3(In6_counter[14]), 
        .IN4(In6_counter[13]), .QN(n703) );
  NAND4X0 U145 ( .IN1(n507), .IN2(n506), .IN3(n505), .IN4(n504), .QN(n711) );
  NOR4X0 U146 ( .IN1(n712), .IN2(In6_counter[6]), .IN3(In6_counter[8]), .IN4(
        In6_counter[7]), .QN(n702) );
  NAND3X0 U147 ( .IN1(n509), .IN2(n508), .IN3(n510), .QN(n712) );
  NAND4X0 U148 ( .IN1(n713), .IN2(n714), .IN3(n715), .IN4(n716), .QN(n675) );
  NOR4X0 U149 ( .IN1(n717), .IN2(In4_counter[24]), .IN3(In4_counter[26]), 
        .IN4(In4_counter[25]), .QN(n716) );
  NAND4X0 U150 ( .IN1(n549), .IN2(n548), .IN3(n547), .IN4(n718), .QN(n717) );
  NAND3X0 U151 ( .IN1(In4_counter[5]), .IN2(In4_counter[4]), .IN3(n719), .QN(
        n718) );
  NAND3X0 U152 ( .IN1(n560), .IN2(n720), .IN3(n561), .QN(n719) );
  NAND2X0 U153 ( .IN1(In4_counter[1]), .IN2(In4_counter[0]), .QN(n720) );
  NOR4X0 U154 ( .IN1(n721), .IN2(In4_counter[18]), .IN3(In4_counter[20]), 
        .IN4(In4_counter[19]), .QN(n715) );
  NAND3X0 U155 ( .IN1(n551), .IN2(n550), .IN3(n552), .QN(n721) );
  NOR4X0 U156 ( .IN1(n722), .IN2(In4_counter[11]), .IN3(In4_counter[13]), 
        .IN4(In4_counter[12]), .QN(n714) );
  NAND4X0 U157 ( .IN1(n556), .IN2(n555), .IN3(n554), .IN4(n553), .QN(n722) );
  NOR4X0 U158 ( .IN1(n723), .IN2(In4_counter[30]), .IN3(In4_counter[7]), .IN4(
        In4_counter[6]), .QN(n713) );
  NAND3X0 U159 ( .IN1(n558), .IN2(n557), .IN3(n559), .QN(n723) );
  NAND4X0 U160 ( .IN1(n724), .IN2(n725), .IN3(n726), .IN4(n727), .QN(n674) );
  NOR4X0 U161 ( .IN1(n728), .IN2(In1_counter[25]), .IN3(In1_counter[27]), 
        .IN4(In1_counter[26]), .QN(n727) );
  NAND4X0 U162 ( .IN1(n516), .IN2(n515), .IN3(n514), .IN4(n729), .QN(n728) );
  NAND3X0 U163 ( .IN1(In1_counter[5]), .IN2(In1_counter[4]), .IN3(n730), .QN(
        n729) );
  NAND3X0 U164 ( .IN1(n527), .IN2(n731), .IN3(n528), .QN(n730) );
  NAND2X0 U165 ( .IN1(In1_counter[1]), .IN2(In1_counter[0]), .QN(n731) );
  NOR4X0 U166 ( .IN1(n732), .IN2(In1_counter[19]), .IN3(In1_counter[21]), 
        .IN4(In1_counter[20]), .QN(n726) );
  NAND3X0 U167 ( .IN1(n518), .IN2(n517), .IN3(n519), .QN(n732) );
  NOR4X0 U168 ( .IN1(n733), .IN2(In1_counter[12]), .IN3(In1_counter[14]), 
        .IN4(In1_counter[13]), .QN(n725) );
  NAND4X0 U169 ( .IN1(n523), .IN2(n522), .IN3(n521), .IN4(n520), .QN(n733) );
  NOR4X0 U170 ( .IN1(n734), .IN2(In1_counter[6]), .IN3(In1_counter[8]), .IN4(
        In1_counter[7]), .QN(n724) );
  NAND3X0 U171 ( .IN1(n525), .IN2(n524), .IN3(n526), .QN(n734) );
  ISOLANDX1 U172 ( .D(N319), .ISO(n629), .Q(N351) );
  ISOLANDX1 U173 ( .D(N318), .ISO(n629), .Q(N350) );
  ISOLANDX1 U174 ( .D(N317), .ISO(n629), .Q(N349) );
  ISOLANDX1 U175 ( .D(N316), .ISO(n629), .Q(N348) );
  ISOLANDX1 U176 ( .D(N315), .ISO(n629), .Q(N347) );
  ISOLANDX1 U177 ( .D(N314), .ISO(n629), .Q(N346) );
  ISOLANDX1 U178 ( .D(N313), .ISO(n629), .Q(N345) );
  ISOLANDX1 U179 ( .D(N312), .ISO(n629), .Q(N344) );
  ISOLANDX1 U180 ( .D(N311), .ISO(n629), .Q(N343) );
  ISOLANDX1 U181 ( .D(N310), .ISO(n629), .Q(N342) );
  ISOLANDX1 U182 ( .D(N309), .ISO(n629), .Q(N341) );
  ISOLANDX1 U183 ( .D(N308), .ISO(n629), .Q(N340) );
  ISOLANDX1 U184 ( .D(N307), .ISO(n629), .Q(N339) );
  ISOLANDX1 U185 ( .D(N306), .ISO(n629), .Q(N338) );
  ISOLANDX1 U186 ( .D(N305), .ISO(n629), .Q(N337) );
  ISOLANDX1 U187 ( .D(N304), .ISO(n629), .Q(N336) );
  ISOLANDX1 U188 ( .D(N303), .ISO(n629), .Q(N335) );
  ISOLANDX1 U189 ( .D(N302), .ISO(n629), .Q(N334) );
  ISOLANDX1 U190 ( .D(N301), .ISO(n629), .Q(N333) );
  ISOLANDX1 U191 ( .D(N300), .ISO(n629), .Q(N332) );
  ISOLANDX1 U192 ( .D(N299), .ISO(n629), .Q(N331) );
  ISOLANDX1 U193 ( .D(N298), .ISO(n629), .Q(N330) );
  ISOLANDX1 U194 ( .D(N297), .ISO(n629), .Q(N329) );
  ISOLANDX1 U195 ( .D(N296), .ISO(n629), .Q(N328) );
  ISOLANDX1 U196 ( .D(N295), .ISO(n629), .Q(N327) );
  ISOLANDX1 U197 ( .D(N294), .ISO(n629), .Q(N326) );
  ISOLANDX1 U198 ( .D(N293), .ISO(n629), .Q(N325) );
  ISOLANDX1 U199 ( .D(N292), .ISO(n629), .Q(N324) );
  ISOLANDX1 U200 ( .D(N291), .ISO(n629), .Q(N323) );
  ISOLANDX1 U201 ( .D(N290), .ISO(n629), .Q(N322) );
  ISOLANDX1 U202 ( .D(N289), .ISO(n629), .Q(N321) );
  ISOLANDX1 U203 ( .D(N288), .ISO(n629), .Q(N320) );
  OA21X1 U204 ( .IN1(n672), .IN2(n735), .IN3(n759), .Q(n629) );
  AND4X1 U205 ( .IN1(n673), .IN2(Clock_counter[2]), .IN3(n736), .IN4(
        Clock_counter[3]), .Q(n735) );
  NOR2X0 U206 ( .IN1(n760), .IN2(n758), .QN(n736) );
  NAND4X0 U207 ( .IN1(n737), .IN2(n738), .IN3(n739), .IN4(n740), .QN(n672) );
  NOR4X0 U208 ( .IN1(n741), .IN2(Clock_counter[12]), .IN3(Clock_counter[10]), 
        .IN4(Clock_counter[11]), .QN(n740) );
  NAND4X0 U209 ( .IN1(n748), .IN2(n747), .IN3(n746), .IN4(n742), .QN(n741) );
  NAND2X0 U210 ( .IN1(n673), .IN2(Clock_counter[4]), .QN(n742) );
  AND2X1 U211 ( .IN1(Clock_counter[5]), .IN2(Clock_counter[6]), .Q(n673) );
  NOR4X0 U212 ( .IN1(n743), .IN2(Clock_counter[18]), .IN3(Clock_counter[16]), 
        .IN4(Clock_counter[17]), .QN(n739) );
  NAND3X0 U213 ( .IN1(n750), .IN2(n749), .IN3(n751), .QN(n743) );
  NOR4X0 U214 ( .IN1(n744), .IN2(Clock_counter[24]), .IN3(Clock_counter[22]), 
        .IN4(Clock_counter[23]), .QN(n738) );
  NAND3X0 U215 ( .IN1(n753), .IN2(n752), .IN3(n754), .QN(n744) );
  NOR4X0 U216 ( .IN1(n745), .IN2(Clock_counter[30]), .IN3(Clock_counter[28]), 
        .IN4(Clock_counter[29]), .QN(n737) );
  NAND3X0 U217 ( .IN1(n756), .IN2(n755), .IN3(n757), .QN(n745) );
endmodule

module s38584 ( CK, g100, g10122, g10306, g10500, g10527, g113, g11349, g11388, 
        g114, g11418, g11447, g115, g116, g11678, g11770, g120, g12184, g12238, 
        g12300, g12350, g12368, g124, g12422, g12470, g125, g126, g127, g12832, 
        g12833, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, 
        g13272, g134, g135, g13865, g13881, g13895, g13906, g13926, g13966, 
        g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, 
        g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, 
        g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, 
        g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, 
        g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, 
        g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, 
        g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, 
        g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, 
        g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, 
        g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, 
        g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g24161, 
        g24162, g24163, g24164, g24165, g24166, g24167, g24168, g24169, g24170, 
        g24171, g24172, g24173, g24174, g24175, g24176, g24177, g24178, g24179, 
        g24180, g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219, 
        g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, 
        g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, 
        g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, 
        g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, 
        g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, 
        g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, 
        g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, 
        g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, 
        g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, 
        g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, 
        g34956, g34972, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, 
        g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, 
        g7243, g7245, g7257, g7260, g73, g7540, g7916, g7946, g8132, g8178, 
        g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, 
        g8398, g84, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, 
        g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, 
        g8920, g90, g9019, g9048, g91, g92, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g99, test_se, test_si1, 
        test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, test_so4, 
        test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, test_si8, 
        test_so8, test_si9, test_so9, test_si10, test_so10, test_si11, 
        test_so11, test_si12, test_so12, test_si13, test_so13, test_si14, 
        test_so14, test_si15, test_so15, test_si16, test_so16, test_si17, 
        test_so17, test_si18, test_so18, test_si19, test_so19, test_si20, 
        test_so20, test_si21, test_so21, test_si22, test_so22, test_si23, 
        test_so23, test_si24, test_so24, test_si25, test_so25, test_si26, 
        test_so26, test_si27, test_so27, test_si28, test_so28, test_si29, 
        test_so29, test_si30, test_so30, test_si31, test_so31, test_si32, 
        test_so32, test_si33, test_so33, test_si34, test_so34, test_si35, 
        test_so35, test_si36, test_so36, test_si37, test_so37, test_si38, 
        test_so38, test_si39, test_so39, test_si40, test_so40, test_si41, 
        test_so41, test_si42, test_so42, test_si43, test_so43, test_si44, 
        test_so44, test_si45, test_so45, test_si46, test_so46, test_si47, 
        test_so47, test_si48, test_so48, test_si49, test_so49, test_si50, 
        test_so50, test_si51, test_so51, test_si52, test_so52, test_si53, 
        test_so53, test_si54, test_so54, test_si55, test_so55, test_si56, 
        test_so56, test_si57, test_so57, test_si58, test_so58, test_si59, 
        test_so59, test_si60, test_so60, test_si61, test_so61, test_si62, 
        test_so62, test_si63, test_so63, test_si64, test_so64, test_si65, 
        test_so65, test_si66, test_so66, test_si67, test_so67, test_si68, 
        test_so68, test_si69, test_so69, test_si70, test_so70, test_si71, 
        test_so71, test_si72, test_so72, test_si73, test_so73, test_si74, 
        test_so74, test_si75, test_so75, test_si76, test_so76, test_si77, 
        test_so77, test_si78, test_so78, test_si79, test_so79, test_si80, 
        test_so80, test_si81, test_so81, test_si82, test_so82, test_si83, 
        test_so83, test_si84, test_so84, test_si85, test_so85, test_si86, 
        test_so86, test_si87, test_so87, test_si88, test_so88, test_si89, 
        test_so89, test_si90, test_so90, test_si91, test_so91, test_si92, 
        test_so92, test_si93, test_so93, test_si94, test_so94, test_si95, 
        test_so95, test_si96, test_so96, test_si97, test_so97, test_si98, 
        test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, g6745, g6746,
         g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, g73, g84, g90,
         g91, g92, g99, test_se, test_si1, test_si2, test_si3, test_si4,
         test_si5, test_si6, test_si7, test_si8, test_si9, test_si10,
         test_si11, test_si12, test_si13, test_si14, test_si15, test_si16,
         test_si17, test_si18, test_si19, test_si20, test_si21, test_si22,
         test_si23, test_si24, test_si25, test_si26, test_si27, test_si28,
         test_si29, test_si30, test_si31, test_si32, test_si33, test_si34,
         test_si35, test_si36, test_si37, test_si38, test_si39, test_si40,
         test_si41, test_si42, test_si43, test_si44, test_si45, test_si46,
         test_si47, test_si48, test_si49, test_si50, test_si51, test_si52,
         test_si53, test_si54, test_si55, test_si56, test_si57, test_si58,
         test_si59, test_si60, test_si61, test_si62, test_si63, test_si64,
         test_si65, test_si66, test_si67, test_si68, test_si69, test_si70,
         test_si71, test_si72, test_si73, test_si74, test_si75, test_si76,
         test_si77, test_si78, test_si79, test_si80, test_si81, test_si82,
         test_si83, test_si84, test_si85, test_si86, test_si87, test_si88,
         test_si89, test_si90, test_si91, test_si92, test_si93, test_si94,
         test_si95, test_si96, test_si97, test_si98, test_si99, test_si100;
  output g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447,
         g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422,
         g12470, g12832, g12833, g12919, g12923, g13039, g13049, g13068,
         g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
         g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
         g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
         g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
         g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
         g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
         g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
         g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
         g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
         g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
         g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
         g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
         g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
         g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164,
         g24165, g24166, g24167, g24168, g24169, g24170, g24171, g24172,
         g24173, g24174, g24175, g24176, g24177, g24178, g24179, g24180,
         g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219,
         g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588,
         g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030,
         g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327,
         g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793,
         g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975,
         g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935,
         g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201,
         g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238,
         g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597,
         g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923,
         g34925, g34927, g34956, g34972, g7243, g7245, g7257, g7260, g7540,
         g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291,
         g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783,
         g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916,
         g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
         g9615, g9617, g9680, g9682, g9741, g9743, g9817, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   g34956, g5057, g33046, g2771, g34441, g1882, g33982, g2299, g34007,
         g4040, g24276, g2547, g30381, g559, g3243, g30405, g452, g25604,
         g3542, g30416, g5232, g30466, g5813, g25736, g34617, g1744, g33974,
         g5909, g30505, g1802, g33554, g3554, g30432, g6219, g33064, g807,
         g34881, g6031, g847, g24216, g24232, g4172, g34733, g4372, g34882,
         g3512, g33026, g31867, g3490, g25668, g24344, g4235, g1600, g33966,
         g1714, g33550, g3155, g30393, g2236, g29248, g4555, g4571, g3698,
         g24274, g1736, g33973, g1968, g30360, g34460, g5607, g30494, g2657,
         g30384, g24340, g490, g29223, g311, g26881, g772, g34252, g5587,
         g30489, g6177, g29301, g6377, g3167, g33022, g5615, g30496, g4567,
         g33043, g29263, g6287, g30533, g1500, g24256, g2563, g34015, g4776,
         g34031, g4593, g34452, g6199, g34646, g2295, g34001, g1384, g25633,
         g1339, g24259, g5180, g33049, g2844, g34609, g1024, g31869, g30490,
         g3598, g30427, g4264, g21894, g767, g33965, g5853, g34645, g2089,
         g33571, g4933, g34267, g4521, g26971, g5507, g34644, g6291, g30534,
         g294, g33535, g30498, g25728, g25743, g3813, g25684, g562, g25613,
         g608, g34438, g1205, g24244, g3909, g30439, g6259, g30541, g5905,
         g30519, g921, g25621, g2955, g34807, g203, g25599, g24235, g4878,
         g34036, g5204, g30476, g3606, g30429, g1926, g32997, g6215, g33063,
         g3586, g30424, g291, g32977, g4674, g34026, g3570, g30420, g33560,
         g676, g29226, g843, g25619, g4332, g34455, g4153, g30457, g6336,
         g33625, g622, g34790, g3506, g30414, g4558, g26966, g3111, g25656,
         g21270, g30390, g939, g34727, g278, g25594, g4492, g26963, g4864,
         g34034, g1036, g33541, g21245, g28093, g1178, g24236, g3239, g30404,
         g718, g28051, g6195, g29303, g1135, g26917, g6395, g33624, g25219,
         g24337, g554, g34911, g496, g33963, g3853, g34627, g5134, g29282,
         g25676, g2485, g33013, g925, g32981, g5555, g30483, g1798, g32994,
         g28070, g2941, g34806, g3905, g30453, g763, g33539, g6255, g30526,
         g4375, g26951, g4871, g34035, g4722, g34636, g590, g32978, g1632,
         g30348, g24336, g3100, g24250, g1437, g29236, g6154, g29298, g1579,
         g5567, g30499, g1752, g33976, g1917, g32996, g744, g30335, g4737,
         g34637, g6267, g30528, g1442, g24251, g30521, g4477, g26960, g24239,
         g4643, g34259, g5264, g30474, g2610, g33016, g5160, g34643, g5933,
         g30510, g1454, g29239, g753, g26897, g1296, g34729, g3151, g34625,
         g34800, g6727, g24353, g3530, g33029, g4104, g33615, g1532, g24253,
         g24281, g33997, g4754, g34263, g1189, g24237, g2287, g33584, g4273,
         g24280, g1389, g26920, g33548, g5835, g29296, g1171, g30338, g4269,
         g21895, g2399, g33588, g4983, g34041, g5611, g30495, g4572, g29279,
         g3143, g25655, g2898, g34795, g3343, g24269, g3235, g30403, g33042,
         g3566, g30419, g34023, g4961, g28090, g4927, g34642, g2259, g30370,
         g2819, g34448, g26946, g5802, g2852, g34610, g417, g24209, g681,
         g28047, g437, g24206, g26891, g5901, g30504, g2886, g34798, g3494,
         g25669, g5511, g30480, g3518, g33027, g1604, g33972, g5092, g25697,
         g4831, g28099, g4382, g26947, g6386, g24350, g479, g24210, g3965,
         g30455, g28084, g2008, g33993, g736, g3933, g30444, g222, g33537,
         g3050, g25650, g1052, g25625, g2122, g30366, g2465, g33593, g5889,
         g30502, g4495, g33036, g25595, g34462, g3179, g33024, g1728, g33552,
         g2433, g34014, g3835, g29273, g6187, g25748, g4917, g34638, g1070,
         g30341, g822, g26899, g914, g30336, g5339, g4164, g26940, g25622,
         g2807, g34447, g4054, g33613, g6191, g25749, g5077, g25704, g5523,
         g33053, g3680, g6637, g30555, g174, g25601, g1682, g33971, g355,
         g26892, g1087, g1105, g26915, g33008, g6307, g30538, g3802, g6159,
         g25750, g2255, g30369, g2815, g34446, g911, g29230, g43, g1748,
         g33975, g5551, g30497, g3558, g30418, g5499, g25721, g34622, g3901,
         g30438, g4888, g34266, g6251, g30540, g1373, g32986, g25648, g157,
         g33960, g2783, g34442, g4281, g3574, g30421, g2112, g33573, g1283,
         g34730, g24205, g4297, g758, g32979, g4639, g34025, g6537, g25763,
         g5543, g30481, g5961, g30517, g6243, g30539, g34880, g24242, g30436,
         g3476, g29265, g1664, g32990, g1246, g24245, g6629, g30553, g246,
         g26907, g4049, g24278, g26955, g2932, g24282, g4575, g29276, g4098,
         g31894, g4498, g33037, g528, g26894, g3139, g25654, g20901, g33962,
         g4584, g34451, g142, g34250, g5831, g29295, g239, g26905, g1216,
         g25629, g2848, g34792, g5022, g25703, g1030, g32983, g13881, g3231,
         g30402, g25757, g1430, g2241, g33999, g1564, g24262, g25729, g6148,
         g9682, g6649, g30558, g110, g225, g26901, g26961, g4504, g33039,
         g5873, g33059, g5037, g31899, g2319, g33007, g5495, g25720, g21891,
         g5208, g30462, g5579, g30487, g5869, g33058, g1589, g24261, g5752,
         g25730, g6279, g30531, g30506, g2975, g34804, g6167, g25747, g2599,
         g33601, g1448, g26922, g2370, g29250, g5164, g30459, g1333, g153,
         g33534, g6549, g30543, g4087, g29275, g34030, g2984, g34980, g3961,
         g30451, g962, g25627, g101, g6625, g30552, g1018, g30337, g24254,
         g4045, g24277, g1467, g29237, g2461, g30378, g33019, g5990, g33623,
         g1256, g29235, g5029, g31902, g6519, g29306, g4169, g1816, g33978,
         g4369, g26970, g4578, g29278, g4459, g34253, g3831, g29272, g2514,
         g33595, g3288, g33610, g33589, g2145, g34605, g1700, g30350, g513,
         g25611, g2841, g5297, g33619, g2763, g34022, g4793, g34033, g952,
         g34726, g1263, g31870, g1950, g33985, g5138, g29283, g2307, g34003,
         g25677, g4664, g34463, g2223, g33006, g5808, g29292, g6645, g30557,
         g2016, g33989, g3873, g33033, g2315, g34005, g2811, g26932, g5957,
         g30516, g2047, g33575, g33032, g5575, g30486, g3752, g25678, g3917,
         g30440, g11447, g1585, g4388, g26949, g6275, g30530, g6311, g30542,
         g1041, g25624, g30383, g2537, g33597, g21292, g34598, g4430, g26957,
         g26967, g4826, g28102, g6239, g30524, g232, g26903, g5268, g30475,
         g6545, g34647, g30377, g1772, g33553, g5052, g31903, g9615, g25715,
         g1890, g33984, g2629, g33602, g572, g28045, g2130, g34603, g4108,
         g33035, g4308, g475, g24208, g990, g31, g24213, g3990, g33614, g33060,
         g1992, g30362, g3171, g33023, g812, g26898, g832, g25618, g5897,
         g30518, g4455, g26959, g2902, g34801, g333, g26884, g168, g25600,
         g26933, g3684, g28066, g3639, g33612, g3338, g24268, g5406, g25716,
         g269, g26906, g401, g24203, g6040, g24346, g441, g24207, g25701,
         g3808, g29269, g9, g34255, g3957, g30450, g4093, g30456, g1760,
         g32991, g24348, g160, g34249, g2279, g30371, g3498, g29268, g586,
         g29224, g2619, g33017, g1183, g30339, g1608, g33967, g8785, g1779,
         g33559, g2652, g29255, g2193, g30368, g2393, g30375, g661, g28052,
         g4950, g28089, g5535, g33055, g2834, g30392, g1361, g30343, g6235,
         g30523, g1146, g24233, g33018, g150, g32976, g1696, g30349, g6555,
         g33067, g26900, g3881, g33034, g6621, g30551, g3470, g25667, g3897,
         g30452, g518, g25612, g538, g34719, g2606, g33607, g1472, g26923,
         g24211, g5188, g33050, g5689, g24341, g405, g24201, g5216, g30463,
         g6494, g4669, g34464, g996, g24243, g4531, g24335, g2860, g34611,
         g4743, g34262, g6593, g30546, g8291, g25591, g4411, g1413, g30347,
         g6641, g30556, g6, g1936, g33562, g55, g504, g25610, g2587, g33015,
         g4480, g31896, g34004, g30428, g5571, g30485, g3578, g30422, g25714,
         g5827, g29294, g3582, g30423, g6271, g30529, g4688, g34028, g2380,
         g33587, g5196, g30460, g3227, g30401, g33990, g17316, g6541, g29309,
         g3203, g30411, g1668, g33546, g4760, g28085, g262, g26904, g1840,
         g33556, g5467, g25722, g460, g25605, g6209, g33062, g20763, g26893,
         g655, g28050, g34626, g2204, g33583, g5256, g30472, g4608, g34454,
         g794, g34850, g4423, g3689, g24272, g5685, g703, g24214, g862, g26909,
         g3247, g30406, g2040, g33569, g8178, g25694, g4146, g34628, g4633,
         g34458, g1157, g24240, g4732, g34634, g25700, g5817, g29293, g2351,
         g33009, g2648, g33603, g6736, g24355, g4944, g34268, g4072, g25691,
         g26890, g3466, g29264, g4116, g28072, g5041, g31900, g4434, g26956,
         g3827, g29271, g6500, g29304, g3133, g29261, g3333, g28063, g979,
         g4681, g34027, g298, g33961, g33604, g1894, g32995, g2988, g34624,
         g3538, g30415, g301, g33536, g26888, g827, g28055, g24238, g2555,
         g33600, g5011, g28105, g199, g34721, g6523, g29307, g30345, g4601,
         g34453, g854, g32980, g1484, g29238, g4922, g34639, g5080, g25695,
         g5863, g33057, g4581, g26969, g2518, g29253, g2567, g34021, g568,
         g26895, g3263, g30413, g6613, g30549, g24347, g6444, g25758, g2965,
         g34808, g5857, g30501, g33969, g890, g34440, g3562, g30433, g21900,
         g1404, g26921, g3817, g29270, g4501, g33038, g31865, g2724, g26926,
         g4704, g28083, g22, g2878, g34797, g5220, g30478, g617, g34724,
         g24212, g316, g26883, g1277, g32985, g6513, g25761, g336, g26886,
         g2882, g34796, g32982, g1906, g33561, g305, g26880, g8, g2799, g26931,
         g4912, g34641, g4157, g34629, g2541, g33598, g2153, g33576, g550,
         g34720, g255, g26902, g29244, g5240, g30468, g1478, g26924, g3863,
         g33031, g1959, g29245, g3480, g29266, g6653, g30559, g2864, g34794,
         g4894, g28087, g3857, g30435, g25609, g1002, g28057, g776, g34439,
         g28, g1236, g4646, g34260, g2476, g33012, g1657, g32989, g2375,
         g34006, g63, g358, g896, g26910, g28043, g3161, g33021, g2384, g29251,
         g12470, g4616, g34456, g4561, g26968, g2024, g33991, g3451, g2795,
         g26930, g613, g34599, g4527, g28082, g1844, g33557, g5937, g30511,
         g33045, g2523, g30379, g24267, g2643, g34020, g1489, g24249, g25592,
         g30382, g5156, g29285, g23683, g25662, g21896, g1955, g33563, g33622,
         g2273, g33582, g4771, g28086, g6098, g25744, g3147, g29262, g3347,
         g24270, g2269, g33581, g191, g2712, g626, g34849, g2729, g28060,
         g5357, g33618, g34038, g4709, g34032, g2927, g34803, g4340, g34459,
         g5929, g30509, g4907, g34640, g4035, g28069, g2946, g21899, g918,
         g31868, g4082, g26938, g25756, g30363, g577, g30334, g1620, g33970,
         g2831, g30391, g667, g25615, g930, g33540, g3937, g30445, g817,
         g25617, g1249, g24247, g837, g24215, g599, g33964, g5475, g25719,
         g29228, g5949, g30514, g6682, g33627, g904, g24231, g2873, g34615,
         g1854, g30356, g5084, g25696, g5603, g30493, g2495, g33594, g2437,
         g34009, g2102, g30365, g2208, g33004, g34018, g4064, g25685, g4899,
         g34040, g2719, g25639, g4785, g34029, g5583, g30488, g781, g34600,
         g6173, g29300, g2917, g34802, g686, g25614, g1252, g28058, g671,
         g29225, g33580, g6283, g30532, g5527, g33054, g4489, g26962, g1974,
         g33564, g1270, g32984, g4966, g34039, g6227, g33065, g3929, g30443,
         g5503, g29291, g24279, g5925, g30508, g1124, g29232, g4955, g34269,
         g5224, g30464, g2012, g33988, g6203, g30522, g5120, g25708, g2389,
         g30374, g4438, g26953, g2429, g34008, g2787, g34444, g34731, g2675,
         g33606, g24334, g4836, g34265, g1199, g30340, g24257, g5547, g30482,
         g2138, g34604, g2338, g33591, g6247, g30525, g2791, g26929, g30448,
         g1291, g34602, g5945, g30513, g5244, g30469, g2759, g33608, g6741,
         g33626, g785, g34725, g1259, g30342, g3484, g29267, g209, g25593,
         g6609, g30548, g5517, g33052, g2449, g34012, g34017, g2715, g24263,
         g936, g26912, g2098, g30364, g4462, g34254, g604, g34251, g6589,
         g30560, g33983, g429, g24204, g1870, g33980, g34631, g1825, g29243,
         g1008, g25623, g4392, g26950, g3546, g30431, g5236, g30467, g1768,
         g30353, g4854, g34467, g3925, g30442, g6509, g29305, g732, g25616,
         g2504, g29252, g4520, g2185, g33003, g37, g34613, g4031, g2070,
         g33570, g4176, g34734, g24275, g4405, g872, g6181, g29302, g24349,
         g4765, g34264, g5563, g30484, g1395, g25634, g1913, g33567, g2331,
         g33585, g6263, g30527, g3945, g30447, g347, g4473, g34256, g1266,
         g25630, g5489, g29290, g29227, g2748, g31872, g5471, g29287, g4540,
         g31897, g6723, g6605, g30562, g34011, g2173, g33996, g21898, g2491,
         g33014, g4849, g34465, g2169, g33995, g30372, g30545, g20654, g30389,
         g2407, g33590, g2868, g34616, g2767, g26927, g1783, g32992, g1312,
         g25631, g5212, g30477, g4245, g34632, g645, g28046, g4291, g20899,
         g26896, g25602, g1129, g26916, g2227, g33578, g2246, g33579, g1830,
         g30354, g3590, g30425, g392, g24200, g1592, g33544, g6505, g25764,
         g1221, g24246, g5921, g30507, g21176, g26889, g30333, g218, g1932,
         g32998, g1624, g32987, g5062, g25702, g5462, g29286, g2689, g34606,
         g6573, g33070, g1677, g29240, g2028, g32999, g2671, g33605, g24255,
         g26945, g1848, g33558, g20557, g25699, g5485, g29289, g2741, g30388,
         g2638, g29254, g4122, g28074, g4322, g34450, g5941, g30512, g2108,
         g33572, g25, g33551, g595, g33538, g2217, g33005, g24248, g2066,
         g33002, g1152, g24234, g5252, g30471, g2165, g34000, g2571, g34016,
         g5176, g33048, g25628, g2827, g26934, g4859, g34468, g424, g24202,
         g1274, g33542, g2803, g34445, g1821, g33555, g2509, g34013, g5073,
         g28091, g26919, g6633, g30554, g5124, g29281, g6303, g30537, g5069,
         g28092, g2994, g34732, g650, g28049, g1636, g33545, g3921, g30441,
         g29247, g6732, g24354, g1306, g25636, g1061, g26914, g3462, g25670,
         g2181, g33998, g956, g25626, g1756, g33977, g5849, g29297, g4112,
         g28071, g30387, g2197, g33577, g33592, g1046, g26913, g482, g28044,
         g4401, g26948, g1514, g30344, g329, g26885, g6565, g33069, g2950,
         g34621, g1345, g28059, g6533, g25762, g4727, g34633, g24352, g1536,
         g26925, g3941, g30446, g370, g25597, g5694, g24342, g1858, g30357,
         g446, g26908, g3219, g30399, g1811, g29242, g6601, g30547, g2441,
         g34010, g1874, g33986, g34257, g6581, g30544, g6597, g30561, g5008,
         g3610, g30430, g2890, g34799, g1978, g33565, g1612, g33968, g112,
         g2856, g34793, g1982, g33566, g30465, g4119, g28073, g6390, g24351,
         g1542, g30346, g4258, g21893, g4818, g5033, g31904, g4717, g34635,
         g1554, g25637, g3849, g29274, g3199, g30396, g25735, g4975, g34037,
         g790, g34791, g5913, g30520, g1902, g30358, g6163, g29299, g4125,
         g4821, g28096, g4939, g28088, g24241, g3207, g30397, g4483, g30409,
         g5142, g29284, g5248, g30470, g2126, g30367, g3694, g24273, g5481,
         g29288, g1964, g30359, g5097, g25698, g3215, g30398, g4427, g26952,
         g2779, g26928, g26954, g1720, g30351, g1367, g31871, g5112, g19,
         g4145, g26939, g2161, g33994, g376, g25596, g2361, g33586, g21901,
         g582, g31866, g2051, g33000, g1193, g26918, g2327, g30373, g907,
         g28056, g947, g34601, g1834, g30355, g3594, g30426, g2999, g34805,
         g2303, g34002, g28053, g723, g29229, g5703, g33620, g546, g34722,
         g2472, g33599, g5953, g30515, g25649, g1740, g33979, g3550, g30417,
         g3845, g25683, g2116, g33574, g30410, g3913, g30454, g34024, g1687,
         g33547, g2681, g30386, g2533, g33596, g324, g26887, g2697, g34607,
         g4417, g31895, g6561, g33068, g1141, g29233, g24258, g30376, g1710,
         g33549, g6527, g29308, g3255, g30408, g1691, g29241, g2936, g34620,
         g5644, g33621, g5152, g25707, g5352, g24339, g2775, g34443, g2922,
         g34619, g29234, g5893, g30503, g6617, g30550, g2060, g33001, g4512,
         g33040, g5599, g30492, g3401, g25664, g4366, g26944, g20652, g34614,
         g3129, g29260, g5170, g33047, g5821, g25733, g6299, g30536, g2079,
         g29246, g4698, g34261, g3703, g33611, g1559, g25638, g34728, g411,
         g29222, g25742, g3953, g30449, g2704, g34608, g6035, g24345, g1300,
         g25635, g4057, g25686, g5200, g30461, g4843, g34466, g5046, g31901,
         g2250, g29249, g26882, g33041, g2453, g33011, g5841, g25734, g2912,
         g34618, g2357, g33010, g164, g31864, g4253, g34630, g5016, g31898,
         g3119, g25653, g1351, g25632, g32988, g4519, g33616, g5115, g29280,
         g3352, g33609, g6657, g30563, g4552, g33044, g3893, g30437, g3211,
         g30412, g5595, g30491, g3614, g30434, g34612, g3125, g29259, g3821,
         g25681, g4141, g25687, g4570, g33617, g5272, g30479, g2735, g29256,
         g728, g28054, g6295, g30535, g2661, g30385, g1988, g30361, g25705,
         g1548, g24260, g3106, g29257, g4659, g34461, g4358, g34258, g1792,
         g32993, g2084, g33992, g3187, g30394, g4311, g34449, g2583, g34019,
         g1094, g29231, g25682, g4284, g21897, g3191, g30395, g4239, g21892,
         g4180, g691, g28048, g534, g34723, g385, g25598, g2004, g33987, g2527,
         g30380, g5456, g26965, g25706, g4507, g30458, g5348, g24338, g3223,
         g30400, g2970, g34623, g5698, g24343, g5260, g30473, g1521, g24252,
         g3522, g33028, g3115, g29258, g3251, g30407, g26958, g34457, g1996,
         g33568, g25663, g4515, g26964, g4300, g34735, g30352, g1379, g33543,
         g24271, g1878, g33981, g5619, g30500, g71, g20049, g29277, g34970,
         g34783, g24266, g28753, g29218, g25689, g34649, g27831, g34978,
         g33894, g18597, g34974, g31521, g34781, g34971, g34977, g25690,
         g25688, g34976, g34657, g34975, g34979, g34843, g24298, DFF_24_n1,
         DFF_150_n1, DFF_178_n1, DFF_206_n1, DFF_228_n1, DFF_348_n1,
         DFF_418_n1, DFF_420_n1, DFF_477_n1, DFF_480_n1, DFF_491_n1,
         DFF_514_n1, DFF_672_n1, DFF_709_n1, DFF_829_n1, DFF_909_n1,
         DFF_944_n1, DFF_961_n1, DFF_992_n1, DFF_1012_n1, DFF_1092_n1,
         DFF_1225_n1, DFF_1234_n1, DFF_1322_n1, DFF_1338_n1, DFF_1381_n1,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1452, n1453, n1454, n1455, n1456, n1457,
         n1461, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1492, n1496,
         n1497, n1498, n1499, n1502, n1503, n1504, n1509, n1510, n1511, n1513,
         n1514, n1516, n1519, n1522, n1523, n1527, n1532, n1534, n1535, n1538,
         n1539, n1540, n1544, n1546, n1548, n1549, n1552, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1570, n1571, n1572, n1573, n1574, n1576, n1577, n1578, g32975, n1581,
         n1582, n1583, n1589, n1590, n1591, n1594, n1599, n1600, n1601, n1602,
         n1604, n1605, n1606, n1607, n1608, n1609, n1611, n1612, n1613, n1621,
         n1622, n1624, n1625, n1634, n1635, n1640, n1641, n1645, n1648, n1650,
         n1655, n1660, n1661, n1666, n1668, n1669, n1670, n1674, n1675, n1676,
         n1678, n1679, n1680, n1681, n1682, n1686, n1692, n1693, n1694, n1695,
         n1696, n1700, n1701, n1702, n1703, n1704, n1705, n1707, n1712, n1713,
         n1715, n1719, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1740,
         n1742, n1743, n1744, n1745, n1747, n1748, n1749, n1751, n1755, n1757,
         n1759, n1761, n1762, n1770, n1775, n1776, n1788, n1790, n1791, n1793,
         n1794, n1795, n1800, n1801, n1802, n1809, n1810, n1816, n1817, n1818,
         n1820, n1821, n1822, n1823, n1824, n1835, n1837, n1840, n1842, n1843,
         n1844, n1845, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1866, n1867, n1869, n1870, n1871,
         n1874, n1877, n1880, n1881, n1882, n1883, n1888, n1890, n1891, n1893,
         g31860, n1903, n1904, n1905, n1907, n1908, n1927, n1928, n1936, n1940,
         n1941, n1942, n1943, n1946, n1952, n1954, n1967, n1968, n1969, n1970,
         n1986, n1987, n1989, g31862, n2004, n2011, n2034, n2035, n2042, n2048,
         n2049, n2063, n2072, g31863, n2075, n2076, n2077, n2101, n2102, n2103,
         n2108, n2119, n2120, n2122, n2123, n2131, n2134, n2135, n2136, n2138,
         n2140, n2172, n2218, n2222, n2223, n2224, n2225, n2226, n2228, n2303,
         n2304, n2305, n2307, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2490, n2492, n2493, n2494, n2496,
         n2497, n2498, n2499, n2500, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2512, n2513, n2514, n2515, n2516, n2518, n2519,
         n2521, n2522, n2523, n2524, n2525, n2527, n2528, n2529, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2540, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3652, n3653, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4875, n4876, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4987, n4988, n4989, n4990, n4992,
         n4993, n4994, n4995, n4997, n4998, n4999, n5000, n5002, n5003, n5004,
         n5005, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5035, n5036,
         n5037, n5038, n5040, n5041, n5042, n5043, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, g34436,
         g34437, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, g30329, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, g23002, g23759,
         g30330, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5896, n5898, n5900, n5902, n5904, n5906, n5908,
         n5910, n5912, n5914, n5916, n5918, n5920, n5922, n5924, n5926, n5928,
         n5930, n5932, n5934, n5936, n5938, n5940, n5942, n5944, n5946, n5948,
         n5950, n5952, n5954, n5956, n5958, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6016, n6018,
         n6021, n6022, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n9236, n9240, n9245, n9247, n9255, n9262, n9265,
         n9267, n9273, n9274, n9276, n9280, n9281, n9294, n9295, n9302, n9303,
         n9306, n9312, n9314, n9322, n9324, n9325, n9327, n9332, n9336, n9340,
         n9348, n9351, n9352, n9357, n9367, g10122_Tj, Tj_Trigger;
  assign g34839 = g34956;
  assign g29217 = g21270;
  assign g29220 = g21245;
  assign test_so10 = g25219;
  assign g31861 = g25219;
  assign g29215 = g20901;
  assign test_so26 = g13881;
  assign test_so92 = g9682;
  assign test_so86 = g11447;
  assign g29221 = g21292;
  assign test_so35 = g9615;
  assign test_so39 = g8785;
  assign test_so42 = g8291;
  assign test_so44 = g17316;
  assign g29211 = g20763;
  assign test_so46 = g8178;
  assign test_so80 = g12470;
  assign g30332 = g23683;
  assign g29219 = g20654;
  assign g29212 = g20899;
  assign g29216 = g21176;
  assign g29213 = g20557;
  assign g29214 = g20652;
  assign test_so100 = g20049;
  assign g29210 = g20049;
  assign g33959 = g28753;
  assign g18881 = g29218;
  assign g33533 = g27831;
  assign g34788 = g33894;
  assign g34435 = g31521;
  assign g26801 = g32975;
  assign g25114 = g31860;
  assign g25259 = g31862;
  assign g25167 = g31863;
  assign g34237 = 1'b1;
  assign g34238 = 1'b1;
  assign g34240 = 1'b1;
  assign g34239 = 1'b1;
  assign g34236 = 1'b1;
  assign g34233 = 1'b1;
  assign g34234 = 1'b1;
  assign g34235 = 1'b1;
  assign g31656 = g34436;
  assign g31665 = g34437;
  assign g34597 = 1'b0;
  assign g33950 = 1'b1;
  assign g33945 = 1'b1;
  assign g32429 = 1'b1;
  assign g34232 = 1'b1;
  assign g33947 = 1'b1;
  assign g33949 = 1'b1;
  assign g33946 = 1'b1;
  assign g33948 = 1'b1;
  assign g32454 = 1'b1;
  assign g25582 = 1'b1;
  assign g25583 = 1'b1;
  assign g25584 = 1'b1;
  assign g25585 = 1'b1;
  assign g25586 = 1'b1;
  assign g25587 = 1'b1;
  assign g25588 = 1'b1;
  assign g25589 = 1'b1;
  assign g25590 = 1'b1;
  assign g24151 = 1'b1;
  assign g23612 = g30329;
  assign g30327 = g23002;
  assign g30331 = g23759;
  assign g23652 = g30330;

  LSDNENX1 U5116 ( .D(g34783), .ENB(n2730), .Q(g34221) );
  LSDNENX1 U5126 ( .D(n4836), .ENB(n4896), .Q(n4895) );
  LSDNENX1 U5127 ( .D(n4837), .ENB(n4921), .Q(n4920) );
  LSDNENX1 U5128 ( .D(n2787), .ENB(n4411), .Q(n5045) );
  LSDNENX1 U5129 ( .D(g559), .ENB(g9048), .Q(n4959) );
  SDFFX1 DFF_0_Q_reg ( .D(g33046), .SI(test_si1), .SE(test_se), .CLK(CK), .Q(
        g5057), .QN(n5615) );
  SDFFX1 DFF_1_Q_reg ( .D(g34441), .SI(g5057), .SE(test_se), .CLK(CK), .Q(
        g2771), .QN(n5544) );
  SDFFX1 DFF_2_Q_reg ( .D(g33982), .SI(g2771), .SE(test_se), .CLK(CK), .Q(
        g1882), .QN(n5854) );
  SDFFX1 DFF_4_Q_reg ( .D(g34007), .SI(g1882), .SE(test_se), .CLK(CK), .Q(
        g2299), .QN() );
  SDFFX1 DFF_5_Q_reg ( .D(g24276), .SI(g2299), .SE(test_se), .CLK(CK), .Q(
        g4040), .QN(n5530) );
  SDFFX1 DFF_6_Q_reg ( .D(g30381), .SI(g4040), .SE(test_se), .CLK(CK), .Q(
        g2547), .QN(n5782) );
  SDFFX1 DFF_7_Q_reg ( .D(g9048), .SI(g2547), .SE(test_se), .CLK(CK), .Q(g559), 
        .QN() );
  SDFFX1 DFF_9_Q_reg ( .D(g30405), .SI(g559), .SE(test_se), .CLK(CK), .Q(g3243), .QN() );
  SDFFX1 DFF_10_Q_reg ( .D(g25604), .SI(g3243), .SE(test_se), .CLK(CK), .Q(
        g452), .QN() );
  SDFFX1 DFF_12_Q_reg ( .D(g30416), .SI(g452), .SE(test_se), .CLK(CK), .Q(
        g3542), .QN() );
  SDFFX1 DFF_13_Q_reg ( .D(g30466), .SI(g3542), .SE(test_se), .CLK(CK), .Q(
        g5232), .QN() );
  SDFFX1 DFF_14_Q_reg ( .D(g25736), .SI(g5232), .SE(test_se), .CLK(CK), .Q(
        g5813), .QN() );
  SDFFX1 DFF_15_Q_reg ( .D(g34617), .SI(g5813), .SE(test_se), .CLK(CK), .Q(
        test_so1), .QN() );
  SDFFX1 DFF_16_Q_reg ( .D(g33974), .SI(test_si2), .SE(test_se), .CLK(CK), .Q(
        g1744), .QN(n5795) );
  SDFFX1 DFF_17_Q_reg ( .D(g30505), .SI(g1744), .SE(test_se), .CLK(CK), .Q(
        g5909), .QN() );
  SDFFX1 DFF_18_Q_reg ( .D(g33554), .SI(g5909), .SE(test_se), .CLK(CK), .Q(
        g1802), .QN(n5536) );
  SDFFX1 DFF_19_Q_reg ( .D(g30432), .SI(g1802), .SE(test_se), .CLK(CK), .Q(
        g3554), .QN() );
  SDFFX1 DFF_20_Q_reg ( .D(g33064), .SI(g3554), .SE(test_se), .CLK(CK), .Q(
        g6219), .QN(n5385) );
  SDFFX1 DFF_21_Q_reg ( .D(g34881), .SI(g6219), .SE(test_se), .CLK(CK), .Q(
        g807), .QN(n5479) );
  SDFFX1 DFF_22_Q_reg ( .D(g17715), .SI(g807), .SE(test_se), .CLK(CK), .Q(
        g6031), .QN() );
  SDFFX1 DFF_23_Q_reg ( .D(g24216), .SI(g6031), .SE(test_se), .CLK(CK), .Q(
        g847), .QN(n5709) );
  SDFFX1 DFF_24_Q_reg ( .D(g24232), .SI(g847), .SE(test_se), .CLK(CK), .Q(
        n9367), .QN(DFF_24_n1) );
  SDFFX1 DFF_25_Q_reg ( .D(g34733), .SI(n9367), .SE(test_se), .CLK(CK), .Q(
        g4172), .QN(n5493) );
  SDFFX1 DFF_26_Q_reg ( .D(g34882), .SI(g4172), .SE(test_se), .CLK(CK), .Q(
        g4372), .QN() );
  SDFFX1 DFF_27_Q_reg ( .D(g33026), .SI(g4372), .SE(test_se), .CLK(CK), .Q(
        g3512), .QN() );
  SDFFX1 DFF_28_Q_reg ( .D(g31867), .SI(g3512), .SE(test_se), .CLK(CK), .Q(
        test_so2), .QN(n5471) );
  SDFFX1 DFF_29_Q_reg ( .D(g25668), .SI(test_si3), .SE(test_se), .CLK(CK), .Q(
        g3490), .QN(n5454) );
  SDFFX1 DFF_30_Q_reg ( .D(g24344), .SI(g3490), .SE(test_se), .CLK(CK), .Q(
        g12350), .QN(n5432) );
  SDFFX1 DFF_31_Q_reg ( .D(g8920), .SI(g12350), .SE(test_se), .CLK(CK), .Q(
        g4235), .QN() );
  SDFFX1 DFF_32_Q_reg ( .D(g33966), .SI(g4235), .SE(test_se), .CLK(CK), .Q(
        g1600), .QN(n5811) );
  SDFFX1 DFF_33_Q_reg ( .D(g33550), .SI(g1600), .SE(test_se), .CLK(CK), .Q(
        g1714), .QN(n5460) );
  SDFFX1 DFF_34_Q_reg ( .D(g16656), .SI(g1714), .SE(test_se), .CLK(CK), .Q(
        g14451), .QN() );
  SDFFX1 DFF_35_Q_reg ( .D(g30393), .SI(g14451), .SE(test_se), .CLK(CK), .Q(
        g3155), .QN(n5366) );
  SDFFX1 DFF_37_Q_reg ( .D(g29248), .SI(g3155), .SE(test_se), .CLK(CK), .Q(
        g2236), .QN() );
  SDFFX1 DFF_38_Q_reg ( .D(g4571), .SI(g2236), .SE(test_se), .CLK(CK), .Q(
        g4555), .QN() );
  SDFFX1 DFF_39_Q_reg ( .D(g24274), .SI(g4555), .SE(test_se), .CLK(CK), .Q(
        g3698), .QN() );
  SDFFX1 DFF_41_Q_reg ( .D(g33973), .SI(g3698), .SE(test_se), .CLK(CK), .Q(
        g1736), .QN(n5817) );
  SDFFX1 DFF_42_Q_reg ( .D(g30360), .SI(g1736), .SE(test_se), .CLK(CK), .Q(
        g1968), .QN(n5664) );
  SDFFX1 DFF_43_Q_reg ( .D(g34460), .SI(g1968), .SE(test_se), .CLK(CK), .Q(
        test_so3), .QN(n5391) );
  SDFFX1 DFF_44_Q_reg ( .D(g30494), .SI(test_si4), .SE(test_se), .CLK(CK), .Q(
        g5607), .QN() );
  SDFFX1 DFF_45_Q_reg ( .D(g30384), .SI(g5607), .SE(test_se), .CLK(CK), .Q(
        g2657), .QN(n5316) );
  SDFFX1 DFF_46_Q_reg ( .D(g24340), .SI(g2657), .SE(test_se), .CLK(CK), .Q(
        g12300), .QN(n5439) );
  SDFFX1 DFF_47_Q_reg ( .D(g29223), .SI(g12300), .SE(test_se), .CLK(CK), .Q(
        g490), .QN(n5708) );
  SDFFX1 DFF_48_Q_reg ( .D(g26881), .SI(g490), .SE(test_se), .CLK(CK), .Q(g311), .QN(n5317) );
  SDFFX1 DFF_50_Q_reg ( .D(g34252), .SI(g311), .SE(test_se), .CLK(CK), .Q(g772), .QN(n5334) );
  SDFFX1 DFF_51_Q_reg ( .D(g30489), .SI(g772), .SE(test_se), .CLK(CK), .Q(
        g5587), .QN() );
  SDFFX1 DFF_52_Q_reg ( .D(g29301), .SI(g5587), .SE(test_se), .CLK(CK), .Q(
        g6177), .QN(n5874) );
  SDFFX1 DFF_53_Q_reg ( .D(g17743), .SI(g6177), .SE(test_se), .CLK(CK), .Q(
        g6377), .QN() );
  SDFFX1 DFF_54_Q_reg ( .D(g33022), .SI(g6377), .SE(test_se), .CLK(CK), .Q(
        g3167), .QN(n5652) );
  SDFFX1 DFF_55_Q_reg ( .D(g30496), .SI(g3167), .SE(test_se), .CLK(CK), .Q(
        g5615), .QN() );
  SDFFX1 DFF_56_Q_reg ( .D(g33043), .SI(g5615), .SE(test_se), .CLK(CK), .Q(
        g4567), .QN() );
  SDFFX1 DFF_58_Q_reg ( .D(g29263), .SI(g4567), .SE(test_se), .CLK(CK), .Q(
        test_so4), .QN(n5746) );
  SDFFX1 DFF_59_Q_reg ( .D(g30533), .SI(test_si5), .SE(test_se), .CLK(CK), .Q(
        g6287), .QN() );
  SDFFX1 DFF_60_Q_reg ( .D(g24256), .SI(g6287), .SE(test_se), .CLK(CK), .Q(
        g1500), .QN(n5302) );
  SDFFX1 DFF_61_Q_reg ( .D(g34015), .SI(g1500), .SE(test_se), .CLK(CK), .Q(
        g2563), .QN(n5816) );
  SDFFX1 DFF_62_Q_reg ( .D(g34031), .SI(g2563), .SE(test_se), .CLK(CK), .Q(
        g4776), .QN(n5707) );
  SDFFX1 DFF_63_Q_reg ( .D(g34452), .SI(g4776), .SE(test_se), .CLK(CK), .Q(
        g4593), .QN(n5303) );
  SDFFX1 DFF_64_Q_reg ( .D(g34646), .SI(g4593), .SE(test_se), .CLK(CK), .Q(
        g6199), .QN(n5644) );
  SDFFX1 DFF_65_Q_reg ( .D(g34001), .SI(g6199), .SE(test_se), .CLK(CK), .Q(
        g2295), .QN(n5815) );
  SDFFX1 DFF_66_Q_reg ( .D(g25633), .SI(g2295), .SE(test_se), .CLK(CK), .Q(
        g1384), .QN() );
  SDFFX1 DFF_67_Q_reg ( .D(g24259), .SI(g1384), .SE(test_se), .CLK(CK), .Q(
        g1339), .QN(n5381) );
  SDFFX1 DFF_68_Q_reg ( .D(g33049), .SI(g1339), .SE(test_se), .CLK(CK), .Q(
        g5180), .QN(n5384) );
  SDFFX1 DFF_69_Q_reg ( .D(g34609), .SI(g5180), .SE(test_se), .CLK(CK), .Q(
        g2844), .QN() );
  SDFFX1 DFF_70_Q_reg ( .D(g31869), .SI(g2844), .SE(test_se), .CLK(CK), .Q(
        g1024), .QN() );
  SDFFX1 DFF_71_Q_reg ( .D(g30490), .SI(g1024), .SE(test_se), .CLK(CK), .Q(
        test_so5), .QN() );
  SDFFX1 DFF_72_Q_reg ( .D(g30427), .SI(test_si6), .SE(test_se), .CLK(CK), .Q(
        g3598), .QN() );
  SDFFX1 DFF_73_Q_reg ( .D(g21894), .SI(g3598), .SE(test_se), .CLK(CK), .Q(
        g4264), .QN(n5823) );
  SDFFX1 DFF_74_Q_reg ( .D(g33965), .SI(g4264), .SE(test_se), .CLK(CK), .Q(
        g767), .QN(n5333) );
  SDFFX1 DFF_75_Q_reg ( .D(g34645), .SI(g767), .SE(test_se), .CLK(CK), .Q(
        g5853), .QN(n5499) );
  SDFFX1 DFF_76_Q_reg ( .D(g16874), .SI(g5853), .SE(test_se), .CLK(CK), .Q(
        g13865), .QN(n5580) );
  SDFFX1 DFF_77_Q_reg ( .D(g33571), .SI(g13865), .SE(test_se), .CLK(CK), .Q(
        g2089), .QN() );
  SDFFX1 DFF_78_Q_reg ( .D(g34267), .SI(g2089), .SE(test_se), .CLK(CK), .Q(
        g4933), .QN(n5878) );
  SDFFX1 DFF_79_Q_reg ( .D(g26971), .SI(g4933), .SE(test_se), .CLK(CK), .Q(
        g4521), .QN(n5752) );
  SDFFX1 DFF_80_Q_reg ( .D(g34644), .SI(g4521), .SE(test_se), .CLK(CK), .Q(
        g5507), .QN(n5643) );
  SDFFX1 DFF_81_Q_reg ( .D(g16627), .SI(g5507), .SE(test_se), .CLK(CK), .Q(
        g16656), .QN() );
  SDFFX1 DFF_82_Q_reg ( .D(g30534), .SI(g16656), .SE(test_se), .CLK(CK), .Q(
        g6291), .QN() );
  SDFFX1 DFF_83_Q_reg ( .D(g33535), .SI(g6291), .SE(test_se), .CLK(CK), .Q(
        g294), .QN(n5680) );
  SDFFX1 DFF_84_Q_reg ( .D(g30498), .SI(g294), .SE(test_se), .CLK(CK), .Q(
        test_so6), .QN() );
  SDFFX1 DFF_85_Q_reg ( .D(g25728), .SI(test_si7), .SE(test_se), .CLK(CK), .Q(
        g9617), .QN(n5722) );
  SDFFX1 DFF_86_Q_reg ( .D(g25743), .SI(g9617), .SE(test_se), .CLK(CK), .Q(
        g9741), .QN() );
  SDFFX1 DFF_87_Q_reg ( .D(g25684), .SI(g9741), .SE(test_se), .CLK(CK), .Q(
        g3813), .QN() );
  SDFFX1 DFF_88_Q_reg ( .D(g25613), .SI(g3813), .SE(test_se), .CLK(CK), .Q(
        g562), .QN() );
  SDFFX1 DFF_89_Q_reg ( .D(g34438), .SI(g562), .SE(test_se), .CLK(CK), .Q(g608), .QN(n5475) );
  SDFFX1 DFF_90_Q_reg ( .D(g24244), .SI(g608), .SE(test_se), .CLK(CK), .Q(
        g1205), .QN(n5547) );
  SDFFX1 DFF_91_Q_reg ( .D(g30439), .SI(g1205), .SE(test_se), .CLK(CK), .Q(
        g3909), .QN() );
  SDFFX1 DFF_92_Q_reg ( .D(g30541), .SI(g3909), .SE(test_se), .CLK(CK), .Q(
        g6259), .QN() );
  SDFFX1 DFF_93_Q_reg ( .D(g30519), .SI(g6259), .SE(test_se), .CLK(CK), .Q(
        g5905), .QN() );
  SDFFX1 DFF_94_Q_reg ( .D(g25621), .SI(g5905), .SE(test_se), .CLK(CK), .Q(
        g921), .QN() );
  SDFFX1 DFF_95_Q_reg ( .D(g34807), .SI(g921), .SE(test_se), .CLK(CK), .Q(
        g2955), .QN() );
  SDFFX1 DFF_96_Q_reg ( .D(g25599), .SI(g2955), .SE(test_se), .CLK(CK), .Q(
        g203), .QN() );
  SDFFX1 DFF_98_Q_reg ( .D(g24235), .SI(g203), .SE(test_se), .CLK(CK), .Q(
        test_so7), .QN() );
  SDFFX1 DFF_99_Q_reg ( .D(g34036), .SI(test_si8), .SE(test_se), .CLK(CK), .Q(
        g4878), .QN(n5283) );
  SDFFX1 DFF_100_Q_reg ( .D(g30476), .SI(g4878), .SE(test_se), .CLK(CK), .Q(
        g5204), .QN() );
  SDFFX1 DFF_101_Q_reg ( .D(g17580), .SI(g5204), .SE(test_se), .CLK(CK), .Q(
        g17604), .QN() );
  SDFFX1 DFF_102_Q_reg ( .D(g30429), .SI(g17604), .SE(test_se), .CLK(CK), .Q(
        g3606), .QN() );
  SDFFX1 DFF_103_Q_reg ( .D(g32997), .SI(g3606), .SE(test_se), .CLK(CK), .Q(
        g1926), .QN(n5510) );
  SDFFX1 DFF_104_Q_reg ( .D(g33063), .SI(g1926), .SE(test_se), .CLK(CK), .Q(
        g6215), .QN(n5651) );
  SDFFX1 DFF_105_Q_reg ( .D(g30424), .SI(g6215), .SE(test_se), .CLK(CK), .Q(
        g3586), .QN() );
  SDFFX1 DFF_106_Q_reg ( .D(g32977), .SI(g3586), .SE(test_se), .CLK(CK), .Q(
        g291), .QN(n5679) );
  SDFFX1 DFF_107_Q_reg ( .D(g34026), .SI(g291), .SE(test_se), .CLK(CK), .Q(
        g4674), .QN(n5440) );
  SDFFX1 DFF_108_Q_reg ( .D(g30420), .SI(g4674), .SE(test_se), .CLK(CK), .Q(
        g3570), .QN() );
  SDFFX1 DFF_109_Q_reg ( .D(g12368), .SI(g3570), .SE(test_se), .CLK(CK), .Q(
        g9048), .QN() );
  SDFFX1 DFF_110_Q_reg ( .D(g17739), .SI(g9048), .SE(test_se), .CLK(CK), .Q(
        g17607), .QN() );
  SDFFX1 DFF_111_Q_reg ( .D(g33560), .SI(g17607), .SE(test_se), .CLK(CK), .Q(
        test_so8), .QN(n5354) );
  SDFFX1 DFF_112_Q_reg ( .D(g29226), .SI(test_si9), .SE(test_se), .CLK(CK), 
        .Q(g676), .QN(n5751) );
  SDFFX1 DFF_113_Q_reg ( .D(g25619), .SI(g676), .SE(test_se), .CLK(CK), .Q(
        g843), .QN() );
  SDFFX1 DFF_115_Q_reg ( .D(g34455), .SI(g843), .SE(test_se), .CLK(CK), .Q(
        g4332), .QN(n5540) );
  SDFFX1 DFF_116_Q_reg ( .D(g30457), .SI(g4332), .SE(test_se), .CLK(CK), .Q(
        g4153), .QN() );
  SDFFX1 DFF_117_Q_reg ( .D(g14694), .SI(g4153), .SE(test_se), .CLK(CK), .Q(
        g17711), .QN() );
  SDFFX1 DFF_118_Q_reg ( .D(g33625), .SI(g17711), .SE(test_se), .CLK(CK), .Q(
        g6336), .QN(n5592) );
  SDFFX1 DFF_119_Q_reg ( .D(g34790), .SI(g6336), .SE(test_se), .CLK(CK), .Q(
        g622), .QN(n5672) );
  SDFFX1 DFF_120_Q_reg ( .D(g30414), .SI(g622), .SE(test_se), .CLK(CK), .Q(
        g3506), .QN(n5576) );
  SDFFX1 DFF_121_Q_reg ( .D(g26966), .SI(g3506), .SE(test_se), .CLK(CK), .Q(
        g4558), .QN() );
  SDFFX1 DFF_123_Q_reg ( .D(g17649), .SI(g4558), .SE(test_se), .CLK(CK), .Q(
        g17685), .QN() );
  SDFFX1 DFF_124_Q_reg ( .D(g25656), .SI(g17685), .SE(test_se), .CLK(CK), .Q(
        g3111), .QN() );
  SDFFX1 DFF_125_Q_reg ( .D(g30390), .SI(g3111), .SE(test_se), .CLK(CK), .Q(
        g21270), .QN() );
  SDFFX1 DFF_126_Q_reg ( .D(g25688), .SI(g21270), .SE(test_se), .CLK(CK), .Q(
        test_so9), .QN() );
  SDFFX1 DFF_127_Q_reg ( .D(g34727), .SI(test_si10), .SE(test_se), .CLK(CK), 
        .Q(g939), .QN(n5415) );
  SDFFX1 DFF_128_Q_reg ( .D(g25594), .SI(g939), .SE(test_se), .CLK(CK), .Q(
        g278), .QN(n5627) );
  SDFFX1 DFF_129_Q_reg ( .D(g26963), .SI(g278), .SE(test_se), .CLK(CK), .Q(
        g4492), .QN() );
  SDFFX1 DFF_130_Q_reg ( .D(g34034), .SI(g4492), .SE(test_se), .CLK(CK), .Q(
        g4864), .QN(n5318) );
  SDFFX1 DFF_131_Q_reg ( .D(g33541), .SI(g4864), .SE(test_se), .CLK(CK), .Q(
        g1036), .QN() );
  SDFFX1 DFF_132_Q_reg ( .D(g28093), .SI(g1036), .SE(test_se), .CLK(CK), .Q(
        g21245), .QN() );
  SDFFX1 DFF_133_Q_reg ( .D(g24236), .SI(g21245), .SE(test_se), .CLK(CK), .Q(
        g1178), .QN() );
  SDFFX1 DFF_134_Q_reg ( .D(g30404), .SI(g1178), .SE(test_se), .CLK(CK), .Q(
        g3239), .QN() );
  SDFFX1 DFF_135_Q_reg ( .D(g28051), .SI(g3239), .SE(test_se), .CLK(CK), .Q(
        g718), .QN() );
  SDFFX1 DFF_136_Q_reg ( .D(g29303), .SI(g718), .SE(test_se), .CLK(CK), .Q(
        g6195), .QN(n5741) );
  SDFFX1 DFF_137_Q_reg ( .D(g26917), .SI(g6195), .SE(test_se), .CLK(CK), .Q(
        g1135), .QN(n5328) );
  SDFFX1 DFF_139_Q_reg ( .D(g33624), .SI(g1135), .SE(test_se), .CLK(CK), .Q(
        g6395), .QN(n5396) );
  SDFFX1 DFF_141_Q_reg ( .D(g24337), .SI(g6395), .SE(test_se), .CLK(CK), .Q(
        g25219), .QN(n5515) );
  SDFFX1 DFF_142_Q_reg ( .D(g34911), .SI(test_si11), .SE(test_se), .CLK(CK), 
        .Q(g554), .QN() );
  SDFFX1 DFF_143_Q_reg ( .D(g33963), .SI(g554), .SE(test_se), .CLK(CK), .Q(
        g496), .QN() );
  SDFFX1 DFF_144_Q_reg ( .D(g34627), .SI(g496), .SE(test_se), .CLK(CK), .Q(
        g3853), .QN(n5641) );
  SDFFX1 DFF_145_Q_reg ( .D(g29282), .SI(g3853), .SE(test_se), .CLK(CK), .Q(
        g5134), .QN(n5807) );
  SDFFX1 DFF_146_Q_reg ( .D(g17320), .SI(g5134), .SE(test_se), .CLK(CK), .Q(
        g17404), .QN() );
  SDFFX1 DFF_147_Q_reg ( .D(g25676), .SI(g17404), .SE(test_se), .CLK(CK), .Q(
        g8344), .QN(n5721) );
  SDFFX1 DFF_148_Q_reg ( .D(g33013), .SI(g8344), .SE(test_se), .CLK(CK), .Q(
        g2485), .QN(n5509) );
  SDFFX1 DFF_149_Q_reg ( .D(g32981), .SI(g2485), .SE(test_se), .CLK(CK), .Q(
        g925), .QN(n5725) );
  SDFFX1 DFF_150_Q_reg ( .D(g34976), .SI(g925), .SE(test_se), .CLK(CK), .Q(
        n9357), .QN(DFF_150_n1) );
  SDFFX1 DFF_151_Q_reg ( .D(g30483), .SI(n9357), .SE(test_se), .CLK(CK), .Q(
        g5555), .QN() );
  SDFFX1 DFF_152_Q_reg ( .D(g14217), .SI(g5555), .SE(test_se), .CLK(CK), .Q(
        g14096), .QN() );
  SDFFX1 DFF_153_Q_reg ( .D(g32994), .SI(g14096), .SE(test_se), .CLK(CK), .Q(
        g1798), .QN(n5833) );
  SDFFX1 DFF_154_Q_reg ( .D(g28070), .SI(g1798), .SE(test_se), .CLK(CK), .Q(
        test_so11), .QN(n5543) );
  SDFFX1 DFF_155_Q_reg ( .D(g34806), .SI(test_si12), .SE(test_se), .CLK(CK), 
        .Q(g2941), .QN() );
  SDFFX1 DFF_156_Q_reg ( .D(g30453), .SI(g2941), .SE(test_se), .CLK(CK), .Q(
        g3905), .QN() );
  SDFFX1 DFF_157_Q_reg ( .D(g33539), .SI(g3905), .SE(test_se), .CLK(CK), .Q(
        g763), .QN(n5332) );
  SDFFX1 DFF_158_Q_reg ( .D(g30526), .SI(g763), .SE(test_se), .CLK(CK), .Q(
        g6255), .QN() );
  SDFFX1 DFF_159_Q_reg ( .D(g26951), .SI(g6255), .SE(test_se), .CLK(CK), .Q(
        g4375), .QN() );
  SDFFX1 DFF_160_Q_reg ( .D(g34035), .SI(g4375), .SE(test_se), .CLK(CK), .Q(
        g4871), .QN(n5443) );
  SDFFX1 DFF_161_Q_reg ( .D(g34636), .SI(g4871), .SE(test_se), .CLK(CK), .Q(
        g4722), .QN(n5345) );
  SDFFX1 DFF_162_Q_reg ( .D(g32978), .SI(g4722), .SE(test_se), .CLK(CK), .Q(
        g590), .QN(n5472) );
  SDFFX1 DFF_163_Q_reg ( .D(g17722), .SI(g590), .SE(test_se), .CLK(CK), .Q(
        g13099), .QN() );
  SDFFX1 DFF_164_Q_reg ( .D(g30348), .SI(g13099), .SE(test_se), .CLK(CK), .Q(
        g1632), .QN(n5836) );
  SDFFX1 DFF_165_Q_reg ( .D(g24336), .SI(g1632), .SE(test_se), .CLK(CK), .Q(
        g12238), .QN(n5438) );
  SDFFX1 DFF_166_Q_reg ( .D(g8215), .SI(g12238), .SE(test_se), .CLK(CK), .Q(
        g3100), .QN() );
  SDFFX1 DFF_167_Q_reg ( .D(g24250), .SI(g3100), .SE(test_se), .CLK(CK), .Q(
        test_so12), .QN(n5617) );
  SDFFX1 DFF_169_Q_reg ( .D(g29236), .SI(test_si13), .SE(test_se), .CLK(CK), 
        .Q(g1437), .QN(n5696) );
  SDFFX1 DFF_170_Q_reg ( .D(g29298), .SI(g1437), .SE(test_se), .CLK(CK), .Q(
        g6154), .QN(n5747) );
  SDFFX1 DFF_171_Q_reg ( .D(g10527), .SI(g6154), .SE(test_se), .CLK(CK), .Q(
        g1579), .QN() );
  SDFFX1 DFF_172_Q_reg ( .D(g30499), .SI(g1579), .SE(test_se), .CLK(CK), .Q(
        g5567), .QN() );
  SDFFX1 DFF_173_Q_reg ( .D(g33976), .SI(g5567), .SE(test_se), .CLK(CK), .Q(
        g1752), .QN(n5797) );
  SDFFX1 DFF_174_Q_reg ( .D(g32996), .SI(g1752), .SE(test_se), .CLK(CK), .Q(
        g1917), .QN() );
  SDFFX1 DFF_175_Q_reg ( .D(g30335), .SI(g1917), .SE(test_se), .CLK(CK), .Q(
        g744), .QN(n5470) );
  SDFFX1 DFF_177_Q_reg ( .D(g34637), .SI(g744), .SE(test_se), .CLK(CK), .Q(
        g4737), .QN(n5867) );
  SDFFX1 DFF_178_Q_reg ( .D(g25694), .SI(g4737), .SE(test_se), .CLK(CK), .Q(
        g8132), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(g30528), .SI(g8132), .SE(test_se), .CLK(CK), .Q(
        g6267), .QN() );
  SDFFX1 DFF_181_Q_reg ( .D(g16775), .SI(g6267), .SE(test_se), .CLK(CK), .Q(
        g16659), .QN() );
  SDFFX1 DFF_182_Q_reg ( .D(g24251), .SI(g16659), .SE(test_se), .CLK(CK), .Q(
        g1442), .QN() );
  SDFFX1 DFF_183_Q_reg ( .D(g30521), .SI(g1442), .SE(test_se), .CLK(CK), .Q(
        test_so13), .QN() );
  SDFFX1 DFF_184_Q_reg ( .D(g26960), .SI(test_si14), .SE(test_se), .CLK(CK), 
        .Q(g4477), .QN(n5849) );
  SDFFX1 DFF_185_Q_reg ( .D(g24239), .SI(g4477), .SE(test_se), .CLK(CK), .Q(
        g10500), .QN() );
  SDFFX1 DFF_186_Q_reg ( .D(g34259), .SI(g10500), .SE(test_se), .CLK(CK), .Q(
        g4643), .QN(n5382) );
  SDFFX1 DFF_187_Q_reg ( .D(g30474), .SI(g4643), .SE(test_se), .CLK(CK), .Q(
        g5264), .QN() );
  SDFFX1 DFF_188_Q_reg ( .D(g12422), .SI(g5264), .SE(test_se), .CLK(CK), .Q(
        g14779), .QN(n5703) );
  SDFFX1 DFF_189_Q_reg ( .D(g33016), .SI(g14779), .SE(test_se), .CLK(CK), .Q(
        g2610), .QN() );
  SDFFX1 DFF_190_Q_reg ( .D(g34643), .SI(g2610), .SE(test_se), .CLK(CK), .Q(
        g5160), .QN(n5498) );
  SDFFX1 DFF_192_Q_reg ( .D(g30510), .SI(g5160), .SE(test_se), .CLK(CK), .Q(
        g5933), .QN() );
  SDFFX1 DFF_193_Q_reg ( .D(g29239), .SI(g5933), .SE(test_se), .CLK(CK), .Q(
        g1454), .QN(n5866) );
  SDFFX1 DFF_194_Q_reg ( .D(g26897), .SI(g1454), .SE(test_se), .CLK(CK), .Q(
        g753), .QN() );
  SDFFX1 DFF_195_Q_reg ( .D(g34729), .SI(g753), .SE(test_se), .CLK(CK), .Q(
        g1296), .QN() );
  SDFFX1 DFF_196_Q_reg ( .D(g34625), .SI(g1296), .SE(test_se), .CLK(CK), .Q(
        g3151), .QN(n5495) );
  SDFFX1 DFF_197_Q_reg ( .D(g34800), .SI(g3151), .SE(test_se), .CLK(CK), .Q(
        test_so14), .QN() );
  SDFFX1 DFF_198_Q_reg ( .D(g24353), .SI(test_si15), .SE(test_se), .CLK(CK), 
        .Q(g6727), .QN(n5531) );
  SDFFX1 DFF_199_Q_reg ( .D(g33029), .SI(g6727), .SE(test_se), .CLK(CK), .Q(
        g3530), .QN(n5569) );
  SDFFX1 DFF_201_Q_reg ( .D(g33615), .SI(g3530), .SE(test_se), .CLK(CK), .Q(
        g4104), .QN() );
  SDFFX1 DFF_202_Q_reg ( .D(g24253), .SI(g4104), .SE(test_se), .CLK(CK), .Q(
        g1532), .QN() );
  SDFFX1 DFF_203_Q_reg ( .D(g24281), .SI(g1532), .SE(test_se), .CLK(CK), .Q(
        g9251), .QN() );
  SDFFX1 DFF_204_Q_reg ( .D(g33997), .SI(g9251), .SE(test_se), .CLK(CK), .Q(
        n9352), .QN(n5688) );
  SDFFX1 DFF_206_Q_reg ( .D(g34971), .SI(n9352), .SE(test_se), .CLK(CK), .Q(
        n9351), .QN(DFF_206_n1) );
  SDFFX1 DFF_207_Q_reg ( .D(g34263), .SI(n9351), .SE(test_se), .CLK(CK), .Q(
        g4754), .QN(n5877) );
  SDFFX1 DFF_208_Q_reg ( .D(g24237), .SI(g4754), .SE(test_se), .CLK(CK), .Q(
        g1189), .QN(n5642) );
  SDFFX1 DFF_209_Q_reg ( .D(g33584), .SI(g1189), .SE(test_se), .CLK(CK), .Q(
        g2287), .QN(n5353) );
  SDFFX1 DFF_210_Q_reg ( .D(g24280), .SI(g2287), .SE(test_se), .CLK(CK), .Q(
        g4273), .QN(n5764) );
  SDFFX1 DFF_211_Q_reg ( .D(g26920), .SI(g4273), .SE(test_se), .CLK(CK), .Q(
        g1389), .QN() );
  SDFFX1 DFF_212_Q_reg ( .D(g33548), .SI(g1389), .SE(test_se), .CLK(CK), .Q(
        test_so15), .QN(n5758) );
  SDFFX1 DFF_213_Q_reg ( .D(g29296), .SI(test_si16), .SE(test_se), .CLK(CK), 
        .Q(g5835), .QN(n5663) );
  SDFFX1 DFF_214_Q_reg ( .D(g30338), .SI(g5835), .SE(test_se), .CLK(CK), .Q(
        g1171), .QN(n5363) );
  SDFFX1 DFF_215_Q_reg ( .D(g21895), .SI(g1171), .SE(test_se), .CLK(CK), .Q(
        g4269), .QN(n5763) );
  SDFFX1 DFF_216_Q_reg ( .D(g33588), .SI(g4269), .SE(test_se), .CLK(CK), .Q(
        g2399), .QN(n5762) );
  SDFFX1 DFF_218_Q_reg ( .D(g34041), .SI(g2399), .SE(test_se), .CLK(CK), .Q(
        g4983), .QN(n5367) );
  SDFFX1 DFF_219_Q_reg ( .D(g30495), .SI(g4983), .SE(test_se), .CLK(CK), .Q(
        g5611), .QN() );
  SDFFX1 DFF_220_Q_reg ( .D(g16744), .SI(g5611), .SE(test_se), .CLK(CK), .Q(
        g16627), .QN() );
  SDFFX1 DFF_221_Q_reg ( .D(g29279), .SI(g16627), .SE(test_se), .CLK(CK), .Q(
        g4572), .QN() );
  SDFFX1 DFF_222_Q_reg ( .D(g25655), .SI(g4572), .SE(test_se), .CLK(CK), .Q(
        g3143), .QN(n5882) );
  SDFFX1 DFF_223_Q_reg ( .D(g34795), .SI(g3143), .SE(test_se), .CLK(CK), .Q(
        g2898), .QN() );
  SDFFX1 DFF_224_Q_reg ( .D(g24269), .SI(g2898), .SE(test_se), .CLK(CK), .Q(
        g3343), .QN() );
  SDFFX1 DFF_225_Q_reg ( .D(g30403), .SI(g3343), .SE(test_se), .CLK(CK), .Q(
        g3235), .QN() );
  SDFFX1 DFF_226_Q_reg ( .D(g33042), .SI(g3235), .SE(test_se), .CLK(CK), .Q(
        test_so16), .QN() );
  SDFFX1 DFF_227_Q_reg ( .D(g30419), .SI(test_si17), .SE(test_se), .CLK(CK), 
        .Q(g3566), .QN() );
  SDFFX1 DFF_228_Q_reg ( .D(g34023), .SI(g3566), .SE(test_se), .CLK(CK), .Q(
        n9348), .QN(DFF_228_n1) );
  SDFFX1 DFF_229_Q_reg ( .D(g28090), .SI(n9348), .SE(test_se), .CLK(CK), .Q(
        g4961), .QN(n5770) );
  SDFFX1 DFF_231_Q_reg ( .D(g34642), .SI(g4961), .SE(test_se), .CLK(CK), .Q(
        g4927), .QN(n5879) );
  SDFFX1 DFF_232_Q_reg ( .D(g30370), .SI(g4927), .SE(test_se), .CLK(CK), .Q(
        g2259), .QN(n5419) );
  SDFFX1 DFF_233_Q_reg ( .D(g34448), .SI(g2259), .SE(test_se), .CLK(CK), .Q(
        g2819), .QN(n5609) );
  SDFFX1 DFF_234_Q_reg ( .D(g26946), .SI(g2819), .SE(test_se), .CLK(CK), .Q(
        g7257), .QN() );
  SDFFX1 DFF_235_Q_reg ( .D(g9617), .SI(g7257), .SE(test_se), .CLK(CK), .Q(
        g5802), .QN() );
  SDFFX1 DFF_236_Q_reg ( .D(g34610), .SI(g5802), .SE(test_se), .CLK(CK), .Q(
        g2852), .QN() );
  SDFFX1 DFF_237_Q_reg ( .D(g24209), .SI(g2852), .SE(test_se), .CLK(CK), .Q(
        g417), .QN(n5358) );
  SDFFX1 DFF_238_Q_reg ( .D(g28047), .SI(g417), .SE(test_se), .CLK(CK), .Q(
        g681), .QN() );
  SDFFX1 DFF_239_Q_reg ( .D(g24206), .SI(g681), .SE(test_se), .CLK(CK), .Q(
        g437), .QN() );
  SDFFX1 DFF_240_Q_reg ( .D(g26891), .SI(g437), .SE(test_se), .CLK(CK), .Q(
        test_so17), .QN(n5825) );
  SDFFX1 DFF_241_Q_reg ( .D(g30504), .SI(test_si18), .SE(test_se), .CLK(CK), 
        .Q(g5901), .QN() );
  SDFFX1 DFF_242_Q_reg ( .D(g34798), .SI(g5901), .SE(test_se), .CLK(CK), .Q(
        g2886), .QN() );
  SDFFX1 DFF_243_Q_reg ( .D(g25669), .SI(g2886), .SE(test_se), .CLK(CK), .Q(
        g3494), .QN(n5889) );
  SDFFX1 DFF_244_Q_reg ( .D(g30480), .SI(g3494), .SE(test_se), .CLK(CK), .Q(
        g5511), .QN(n5575) );
  SDFFX1 DFF_245_Q_reg ( .D(g33027), .SI(g5511), .SE(test_se), .CLK(CK), .Q(
        g3518), .QN(n5645) );
  SDFFX1 DFF_246_Q_reg ( .D(g33972), .SI(g3518), .SE(test_se), .CLK(CK), .Q(
        g1604), .QN() );
  SDFFX1 DFF_248_Q_reg ( .D(g25697), .SI(g1604), .SE(test_se), .CLK(CK), .Q(
        g5092), .QN() );
  SDFFX1 DFF_249_Q_reg ( .D(g28099), .SI(g5092), .SE(test_se), .CLK(CK), .Q(
        g4831), .QN() );
  SDFFX1 DFF_250_Q_reg ( .D(g26947), .SI(g4831), .SE(test_se), .CLK(CK), .Q(
        g4382), .QN(n5714) );
  SDFFX1 DFF_251_Q_reg ( .D(g24350), .SI(g4382), .SE(test_se), .CLK(CK), .Q(
        g6386), .QN() );
  SDFFX1 DFF_252_Q_reg ( .D(g24210), .SI(g6386), .SE(test_se), .CLK(CK), .Q(
        g479), .QN() );
  SDFFX1 DFF_253_Q_reg ( .D(g30455), .SI(g479), .SE(test_se), .CLK(CK), .Q(
        g3965), .QN() );
  SDFFX1 DFF_254_Q_reg ( .D(g28084), .SI(g3965), .SE(test_se), .CLK(CK), .Q(
        test_so18), .QN(n5773) );
  SDFFX1 DFF_255_Q_reg ( .D(g33993), .SI(test_si19), .SE(test_se), .CLK(CK), 
        .Q(g2008), .QN() );
  SDFFX1 DFF_256_Q_reg ( .D(g11678), .SI(g2008), .SE(test_se), .CLK(CK), .Q(
        g736), .QN() );
  SDFFX1 DFF_257_Q_reg ( .D(g30444), .SI(g736), .SE(test_se), .CLK(CK), .Q(
        g3933), .QN() );
  SDFFX1 DFF_258_Q_reg ( .D(g33537), .SI(g3933), .SE(test_se), .CLK(CK), .Q(
        g222), .QN() );
  SDFFX1 DFF_259_Q_reg ( .D(g25650), .SI(g222), .SE(test_se), .CLK(CK), .Q(
        g3050), .QN(n5998) );
  SDFFX1 DFF_261_Q_reg ( .D(g25625), .SI(g3050), .SE(test_se), .CLK(CK), .Q(
        g1052), .QN() );
  SDFFX1 DFF_263_Q_reg ( .D(g17711), .SI(g1052), .SE(test_se), .CLK(CK), .Q(
        g17580), .QN() );
  SDFFX1 DFF_264_Q_reg ( .D(g30366), .SI(g17580), .SE(test_se), .CLK(CK), .Q(
        g2122), .QN(n5784) );
  SDFFX1 DFF_265_Q_reg ( .D(g33593), .SI(g2122), .SE(test_se), .CLK(CK), .Q(
        g2465), .QN(n5523) );
  SDFFX1 DFF_267_Q_reg ( .D(g30502), .SI(g2465), .SE(test_se), .CLK(CK), .Q(
        g5889), .QN() );
  SDFFX1 DFF_268_Q_reg ( .D(g33036), .SI(g5889), .SE(test_se), .CLK(CK), .Q(
        g4495), .QN() );
  SDFFX1 DFF_269_Q_reg ( .D(g25595), .SI(g4495), .SE(test_se), .CLK(CK), .Q(
        g8719), .QN() );
  SDFFX1 DFF_270_Q_reg ( .D(g34462), .SI(g8719), .SE(test_se), .CLK(CK), .Q(
        test_so19), .QN() );
  SDFFX1 DFF_271_Q_reg ( .D(g33024), .SI(test_si20), .SE(test_se), .CLK(CK), 
        .Q(g3179), .QN(n5390) );
  SDFFX1 DFF_272_Q_reg ( .D(g33552), .SI(g3179), .SE(test_se), .CLK(CK), .Q(
        g1728), .QN(n5352) );
  SDFFX1 DFF_273_Q_reg ( .D(g34014), .SI(g1728), .SE(test_se), .CLK(CK), .Q(
        g2433), .QN() );
  SDFFX1 DFF_274_Q_reg ( .D(g29273), .SI(g2433), .SE(test_se), .CLK(CK), .Q(
        g3835), .QN(n5662) );
  SDFFX1 DFF_275_Q_reg ( .D(g25748), .SI(g3835), .SE(test_se), .CLK(CK), .Q(
        g6187), .QN(n5453) );
  SDFFX1 DFF_276_Q_reg ( .D(g34638), .SI(g6187), .SE(test_se), .CLK(CK), .Q(
        g4917), .QN(n5408) );
  SDFFX1 DFF_277_Q_reg ( .D(g30341), .SI(g4917), .SE(test_se), .CLK(CK), .Q(
        g1070), .QN() );
  SDFFX1 DFF_278_Q_reg ( .D(g26899), .SI(g1070), .SE(test_se), .CLK(CK), .Q(
        g822), .QN(n5422) );
  SDFFX1 DFF_279_Q_reg ( .D(g14673), .SI(g822), .SE(test_se), .CLK(CK), .Q(
        g17715), .QN() );
  SDFFX1 DFF_280_Q_reg ( .D(g30336), .SI(g17715), .SE(test_se), .CLK(CK), .Q(
        g914), .QN(n5560) );
  SDFFX1 DFF_281_Q_reg ( .D(g17639), .SI(g914), .SE(test_se), .CLK(CK), .Q(
        g5339), .QN() );
  SDFFX1 DFF_282_Q_reg ( .D(g26940), .SI(g5339), .SE(test_se), .CLK(CK), .Q(
        g4164), .QN() );
  SDFFX1 DFF_283_Q_reg ( .D(g25622), .SI(g4164), .SE(test_se), .CLK(CK), .Q(
        test_so20), .QN(n5467) );
  SDFFX1 DFF_284_Q_reg ( .D(g34447), .SI(test_si21), .SE(test_se), .CLK(CK), 
        .Q(g2807), .QN(n5379) );
  SDFFX1 DFF_286_Q_reg ( .D(g33613), .SI(g2807), .SE(test_se), .CLK(CK), .Q(
        g4054), .QN(n5395) );
  SDFFX1 DFF_287_Q_reg ( .D(g25749), .SI(g4054), .SE(test_se), .CLK(CK), .Q(
        g6191), .QN(n5888) );
  SDFFX1 DFF_288_Q_reg ( .D(g25704), .SI(g6191), .SE(test_se), .CLK(CK), .Q(
        g5077), .QN(n5455) );
  SDFFX1 DFF_289_Q_reg ( .D(g33053), .SI(g5077), .SE(test_se), .CLK(CK), .Q(
        g5523), .QN(n5647) );
  SDFFX1 DFF_290_Q_reg ( .D(g16722), .SI(g5523), .SE(test_se), .CLK(CK), .Q(
        g3680), .QN() );
  SDFFX1 DFF_291_Q_reg ( .D(g30555), .SI(g3680), .SE(test_se), .CLK(CK), .Q(
        g6637), .QN() );
  SDFFX1 DFF_292_Q_reg ( .D(g25601), .SI(g6637), .SE(test_se), .CLK(CK), .Q(
        g174), .QN(n5402) );
  SDFFX1 DFF_293_Q_reg ( .D(g33971), .SI(g174), .SE(test_se), .CLK(CK), .Q(
        g1682), .QN() );
  SDFFX1 DFF_294_Q_reg ( .D(g26892), .SI(g1682), .SE(test_se), .CLK(CK), .Q(
        g355), .QN() );
  SDFFX1 DFF_295_Q_reg ( .D(g17400), .SI(g355), .SE(test_se), .CLK(CK), .Q(
        g1087), .QN() );
  SDFFX1 DFF_296_Q_reg ( .D(g26915), .SI(g1087), .SE(test_se), .CLK(CK), .Q(
        g1105), .QN(n5478) );
  SDFFX1 DFF_297_Q_reg ( .D(g33008), .SI(g1105), .SE(test_se), .CLK(CK), .Q(
        test_so21), .QN() );
  SDFFX1 DFF_298_Q_reg ( .D(g30538), .SI(test_si22), .SE(test_se), .CLK(CK), 
        .Q(g6307), .QN() );
  SDFFX1 DFF_299_Q_reg ( .D(g8344), .SI(g6307), .SE(test_se), .CLK(CK), .Q(
        g3802), .QN() );
  SDFFX1 DFF_300_Q_reg ( .D(g25750), .SI(g3802), .SE(test_se), .CLK(CK), .Q(
        g6159), .QN() );
  SDFFX1 DFF_301_Q_reg ( .D(g30369), .SI(g6159), .SE(test_se), .CLK(CK), .Q(
        g2255), .QN(n5414) );
  SDFFX1 DFF_302_Q_reg ( .D(g34446), .SI(g2255), .SE(test_se), .CLK(CK), .Q(
        g2815), .QN(n5404) );
  SDFFX1 DFF_303_Q_reg ( .D(g29230), .SI(g2815), .SE(test_se), .CLK(CK), .Q(
        g911), .QN(n5559) );
  SDFFX1 DFF_304_Q_reg ( .D(n1473), .SI(g911), .SE(test_se), .CLK(CK), .Q(g43), 
        .QN() );
  SDFFX1 DFF_305_Q_reg ( .D(g13966), .SI(g43), .SE(test_se), .CLK(CK), .Q(
        g16775), .QN() );
  SDFFX1 DFF_306_Q_reg ( .D(g33975), .SI(g16775), .SE(test_se), .CLK(CK), .Q(
        g1748), .QN(n5853) );
  SDFFX1 DFF_307_Q_reg ( .D(g30497), .SI(g1748), .SE(test_se), .CLK(CK), .Q(
        g5551), .QN() );
  SDFFX1 DFF_309_Q_reg ( .D(g30418), .SI(g5551), .SE(test_se), .CLK(CK), .Q(
        g3558), .QN() );
  SDFFX1 DFF_310_Q_reg ( .D(g25721), .SI(g3558), .SE(test_se), .CLK(CK), .Q(
        g5499), .QN(n5885) );
  SDFFX1 DFF_311_Q_reg ( .D(g34622), .SI(g5499), .SE(test_se), .CLK(CK), .Q(
        test_so22), .QN() );
  SDFFX1 DFF_312_Q_reg ( .D(g30438), .SI(test_si23), .SE(test_se), .CLK(CK), 
        .Q(g3901), .QN() );
  SDFFX1 DFF_313_Q_reg ( .D(g34266), .SI(g3901), .SE(test_se), .CLK(CK), .Q(
        g4888), .QN(n5863) );
  SDFFX1 DFF_314_Q_reg ( .D(g30540), .SI(g4888), .SE(test_se), .CLK(CK), .Q(
        g6251), .QN() );
  SDFFX1 DFF_315_Q_reg ( .D(g17760), .SI(g6251), .SE(test_se), .CLK(CK), .Q(
        g17649), .QN() );
  SDFFX1 DFF_316_Q_reg ( .D(g32986), .SI(g17649), .SE(test_se), .CLK(CK), .Q(
        g1373), .QN() );
  SDFFX1 DFF_317_Q_reg ( .D(g25648), .SI(g1373), .SE(test_se), .CLK(CK), .Q(
        g8215), .QN(n5723) );
  SDFFX1 DFF_318_Q_reg ( .D(g33960), .SI(g8215), .SE(test_se), .CLK(CK), .Q(
        g157), .QN(n5678) );
  SDFFX1 DFF_319_Q_reg ( .D(g34442), .SI(g157), .SE(test_se), .CLK(CK), .Q(
        g2783), .QN(n5403) );
  SDFFX1 DFF_320_Q_reg ( .D(g8839), .SI(g2783), .SE(test_se), .CLK(CK), .Q(
        g4281), .QN() );
  SDFFX1 DFF_321_Q_reg ( .D(g30421), .SI(g4281), .SE(test_se), .CLK(CK), .Q(
        g3574), .QN() );
  SDFFX1 DFF_322_Q_reg ( .D(g33573), .SI(g3574), .SE(test_se), .CLK(CK), .Q(
        g2112), .QN(n5848) );
  SDFFX1 DFF_323_Q_reg ( .D(g34730), .SI(g2112), .SE(test_se), .CLK(CK), .Q(
        g1283), .QN(n5635) );
  SDFFX1 DFF_324_Q_reg ( .D(g24205), .SI(g1283), .SE(test_se), .CLK(CK), .Q(
        test_so23), .QN() );
  SDFFX1 DFF_325_Q_reg ( .D(g10122_Tj), .SI(test_si24), .SE(test_se), .CLK(CK), 
        .Q(g4297), .QN() );
  SDFFX1 DFF_326_Q_reg ( .D(g12350), .SI(g4297), .SE(test_se), .CLK(CK), .Q(
        g14738), .QN(n5698) );
  SDFFX1 DFF_327_Q_reg ( .D(g19357), .SI(g14738), .SE(test_se), .CLK(CK), .Q(
        g13272), .QN() );
  SDFFX1 DFF_328_Q_reg ( .D(g32979), .SI(g13272), .SE(test_se), .CLK(CK), .Q(
        g758), .QN(n5331) );
  SDFFX1 DFF_331_Q_reg ( .D(g34025), .SI(g758), .SE(test_se), .CLK(CK), .Q(
        g4639), .QN(n5727) );
  SDFFX1 DFF_332_Q_reg ( .D(g25763), .SI(g4639), .SE(test_se), .CLK(CK), .Q(
        g6537), .QN(n5884) );
  SDFFX1 DFF_333_Q_reg ( .D(g30481), .SI(g6537), .SE(test_se), .CLK(CK), .Q(
        g5543), .QN() );
  SDFFX1 DFF_334_Q_reg ( .D(n6024), .SI(g5543), .SE(test_se), .CLK(CK), .Q(
        g8475), .QN() );
  SDFFX1 DFF_336_Q_reg ( .D(g30517), .SI(g8475), .SE(test_se), .CLK(CK), .Q(
        g5961), .QN() );
  SDFFX1 DFF_337_Q_reg ( .D(g30539), .SI(g5961), .SE(test_se), .CLK(CK), .Q(
        g6243), .QN() );
  SDFFX1 DFF_338_Q_reg ( .D(g34880), .SI(g6243), .SE(test_se), .CLK(CK), .Q(
        n9340), .QN(n5338) );
  SDFFX1 DFF_339_Q_reg ( .D(g24242), .SI(n9340), .SE(test_se), .CLK(CK), .Q(
        g12919), .QN(n5654) );
  SDFFX1 DFF_340_Q_reg ( .D(g30436), .SI(g12919), .SE(test_se), .CLK(CK), .Q(
        test_so24), .QN() );
  SDFFX1 DFF_341_Q_reg ( .D(g29265), .SI(test_si25), .SE(test_se), .CLK(CK), 
        .Q(g3476), .QN(n5786) );
  SDFFX1 DFF_342_Q_reg ( .D(g32990), .SI(g3476), .SE(test_se), .CLK(CK), .Q(
        g1664), .QN(n5407) );
  SDFFX1 DFF_343_Q_reg ( .D(g24245), .SI(g1664), .SE(test_se), .CLK(CK), .Q(
        g1246), .QN(n5756) );
  SDFFX1 DFF_345_Q_reg ( .D(g30553), .SI(g1246), .SE(test_se), .CLK(CK), .Q(
        g6629), .QN() );
  SDFFX1 DFF_346_Q_reg ( .D(g26907), .SI(g6629), .SE(test_se), .CLK(CK), .Q(
        g246), .QN(n6008) );
  SDFFX1 DFF_347_Q_reg ( .D(g24278), .SI(g246), .SE(test_se), .CLK(CK), .Q(
        g4049), .QN() );
  SDFFX1 DFF_348_Q_reg ( .D(g26955), .SI(g4049), .SE(test_se), .CLK(CK), .Q(
        g7260), .QN(DFF_348_n1) );
  SDFFX1 DFF_349_Q_reg ( .D(g24282), .SI(g7260), .SE(test_se), .CLK(CK), .Q(
        g2932), .QN() );
  SDFFX1 DFF_350_Q_reg ( .D(g29276), .SI(g2932), .SE(test_se), .CLK(CK), .Q(
        g4575), .QN() );
  SDFFX1 DFF_351_Q_reg ( .D(g31894), .SI(g4575), .SE(test_se), .CLK(CK), .Q(
        g4098), .QN(n5350) );
  SDFFX1 DFF_352_Q_reg ( .D(g33037), .SI(g4098), .SE(test_se), .CLK(CK), .Q(
        g4498), .QN() );
  SDFFX1 DFF_353_Q_reg ( .D(g26894), .SI(g4498), .SE(test_se), .CLK(CK), .Q(
        g528), .QN(n5327) );
  SDFFX1 DFF_355_Q_reg ( .D(g34977), .SI(g528), .SE(test_se), .CLK(CK), .Q(
        test_so25), .QN(n5477) );
  SDFFX1 DFF_356_Q_reg ( .D(g25654), .SI(test_si26), .SE(test_se), .CLK(CK), 
        .Q(g3139), .QN(n5447) );
  SDFFX1 DFF_357_Q_reg ( .D(g33962), .SI(g3139), .SE(test_se), .CLK(CK), .Q(
        g20901), .QN() );
  SDFFX1 DFF_358_Q_reg ( .D(g34451), .SI(g20901), .SE(test_se), .CLK(CK), .Q(
        g4584), .QN(n5539) );
  SDFFX1 DFF_359_Q_reg ( .D(g34250), .SI(g4584), .SE(test_se), .CLK(CK), .Q(
        g142), .QN(n5724) );
  SDFFX1 DFF_360_Q_reg ( .D(g14597), .SI(g142), .SE(test_se), .CLK(CK), .Q(
        g17639), .QN() );
  SDFFX1 DFF_361_Q_reg ( .D(g29295), .SI(g17639), .SE(test_se), .CLK(CK), .Q(
        g5831), .QN(n5873) );
  SDFFX1 DFF_362_Q_reg ( .D(g26905), .SI(g5831), .SE(test_se), .CLK(CK), .Q(
        g239), .QN() );
  SDFFX1 DFF_363_Q_reg ( .D(g25629), .SI(g239), .SE(test_se), .CLK(CK), .Q(
        g1216), .QN(n5442) );
  SDFFX1 DFF_364_Q_reg ( .D(g34792), .SI(g1216), .SE(test_se), .CLK(CK), .Q(
        g2848), .QN() );
  SDFFX1 DFF_366_Q_reg ( .D(g25703), .SI(g2848), .SE(test_se), .CLK(CK), .Q(
        g5022), .QN() );
  SDFFX1 DFF_367_Q_reg ( .D(g14518), .SI(g5022), .SE(test_se), .CLK(CK), .Q(
        g16955), .QN() );
  SDFFX1 DFF_368_Q_reg ( .D(g32983), .SI(g16955), .SE(test_se), .CLK(CK), .Q(
        g1030), .QN() );
  SDFFX1 DFF_369_Q_reg ( .D(g16924), .SI(g1030), .SE(test_se), .CLK(CK), .Q(
        g13881), .QN(n5585) );
  SDFFX1 DFF_370_Q_reg ( .D(g30402), .SI(test_si27), .SE(test_se), .CLK(CK), 
        .Q(g3231), .QN() );
  SDFFX1 DFF_371_Q_reg ( .D(g25757), .SI(g3231), .SE(test_se), .CLK(CK), .Q(
        g9817), .QN() );
  SDFFX1 DFF_372_Q_reg ( .D(g17423), .SI(g9817), .SE(test_se), .CLK(CK), .Q(
        g1430), .QN() );
  SDFFX1 DFF_373_Q_reg ( .D(g7245), .SI(g1430), .SE(test_se), .CLK(CK), .Q(
        n9336), .QN(n5819) );
  SDFFX1 DFF_374_Q_reg ( .D(g33999), .SI(n9336), .SE(test_se), .CLK(CK), .Q(
        g2241), .QN() );
  SDFFX1 DFF_375_Q_reg ( .D(g24262), .SI(g2241), .SE(test_se), .CLK(CK), .Q(
        g1564), .QN() );
  SDFFX1 DFF_376_Q_reg ( .D(g25729), .SI(g1564), .SE(test_se), .CLK(CK), .Q(
        g9680), .QN() );
  SDFFX1 DFF_377_Q_reg ( .D(g9682), .SI(g9680), .SE(test_se), .CLK(CK), .Q(
        g6148), .QN() );
  SDFFX1 DFF_378_Q_reg ( .D(g30558), .SI(g6148), .SE(test_se), .CLK(CK), .Q(
        g6649), .QN() );
  SDFFX1 DFF_379_Q_reg ( .D(g34781), .SI(g6649), .SE(test_se), .CLK(CK), .Q(
        g110), .QN() );
  SDFFX1 DFF_380_Q_reg ( .D(g14125), .SI(g110), .SE(test_se), .CLK(CK), .Q(
        g14147), .QN() );
  SDFFX1 DFF_382_Q_reg ( .D(g26901), .SI(g14147), .SE(test_se), .CLK(CK), .Q(
        g225), .QN(n5597) );
  SDFFX1 DFF_383_Q_reg ( .D(g26961), .SI(g225), .SE(test_se), .CLK(CK), .Q(
        test_so27), .QN() );
  SDFFX1 DFF_384_Q_reg ( .D(g33039), .SI(test_si28), .SE(test_se), .CLK(CK), 
        .Q(g4504), .QN() );
  SDFFX1 DFF_385_Q_reg ( .D(g33059), .SI(g4504), .SE(test_se), .CLK(CK), .Q(
        g5873), .QN(n5388) );
  SDFFX1 DFF_386_Q_reg ( .D(g31899), .SI(g5873), .SE(test_se), .CLK(CK), .Q(
        g5037), .QN(n5611) );
  SDFFX1 DFF_387_Q_reg ( .D(g33007), .SI(g5037), .SE(test_se), .CLK(CK), .Q(
        g2319), .QN(n5375) );
  SDFFX1 DFF_388_Q_reg ( .D(g25720), .SI(g2319), .SE(test_se), .CLK(CK), .Q(
        g5495), .QN(n5446) );
  SDFFX1 DFF_389_Q_reg ( .D(g21891), .SI(g5495), .SE(test_se), .CLK(CK), .Q(
        g11770), .QN() );
  SDFFX1 DFF_390_Q_reg ( .D(g30462), .SI(g11770), .SE(test_se), .CLK(CK), .Q(
        g5208), .QN() );
  SDFFX1 DFF_392_Q_reg ( .D(g30487), .SI(g5208), .SE(test_se), .CLK(CK), .Q(
        g5579), .QN() );
  SDFFX1 DFF_393_Q_reg ( .D(g33058), .SI(g5579), .SE(test_se), .CLK(CK), .Q(
        g5869), .QN(n5649) );
  SDFFX1 DFF_395_Q_reg ( .D(g24261), .SI(g5869), .SE(test_se), .CLK(CK), .Q(
        g1589), .QN(n5755) );
  SDFFX1 DFF_396_Q_reg ( .D(g25730), .SI(g1589), .SE(test_se), .CLK(CK), .Q(
        g5752), .QN(n5996) );
  SDFFX1 DFF_397_Q_reg ( .D(g30531), .SI(g5752), .SE(test_se), .CLK(CK), .Q(
        g6279), .QN() );
  SDFFX1 DFF_398_Q_reg ( .D(g30506), .SI(g6279), .SE(test_se), .CLK(CK), .Q(
        test_so28), .QN() );
  SDFFX1 DFF_399_Q_reg ( .D(g34804), .SI(test_si29), .SE(test_se), .CLK(CK), 
        .Q(g2975), .QN(n5750) );
  SDFFX1 DFF_400_Q_reg ( .D(g25747), .SI(g2975), .SE(test_se), .CLK(CK), .Q(
        g6167), .QN(n5430) );
  SDFFX1 DFF_401_Q_reg ( .D(g11418), .SI(g6167), .SE(test_se), .CLK(CK), .Q(
        g13966), .QN(n5701) );
  SDFFX1 DFF_402_Q_reg ( .D(g33601), .SI(g13966), .SE(test_se), .CLK(CK), .Q(
        g2599), .QN(n5524) );
  SDFFX1 DFF_403_Q_reg ( .D(g26922), .SI(g2599), .SE(test_se), .CLK(CK), .Q(
        g1448), .QN(n5343) );
  SDFFX1 DFF_404_Q_reg ( .D(g14096), .SI(g1448), .SE(test_se), .CLK(CK), .Q(
        g14125), .QN() );
  SDFFX1 DFF_406_Q_reg ( .D(g29250), .SI(g14125), .SE(test_se), .CLK(CK), .Q(
        g2370), .QN() );
  SDFFX1 DFF_407_Q_reg ( .D(g30459), .SI(g2370), .SE(test_se), .CLK(CK), .Q(
        g5164), .QN(n5570) );
  SDFFX1 DFF_408_Q_reg ( .D(g8475), .SI(g5164), .SE(test_se), .CLK(CK), .Q(
        g1333), .QN(n5616) );
  SDFFX1 DFF_409_Q_reg ( .D(g33534), .SI(g1333), .SE(test_se), .CLK(CK), .Q(
        g153), .QN(n5677) );
  SDFFX1 DFF_410_Q_reg ( .D(g30543), .SI(g153), .SE(test_se), .CLK(CK), .Q(
        g6549), .QN(n5571) );
  SDFFX1 DFF_411_Q_reg ( .D(g29275), .SI(g6549), .SE(test_se), .CLK(CK), .Q(
        g4087), .QN(n5480) );
  SDFFX1 DFF_412_Q_reg ( .D(g34030), .SI(g4087), .SE(test_se), .CLK(CK), .Q(
        test_so29), .QN(n5285) );
  SDFFX1 DFF_413_Q_reg ( .D(g34980), .SI(test_si30), .SE(test_se), .CLK(CK), 
        .Q(g2984), .QN(n5842) );
  SDFFX1 DFF_414_Q_reg ( .D(g30451), .SI(g2984), .SE(test_se), .CLK(CK), .Q(
        g3961), .QN() );
  SDFFX1 DFF_416_Q_reg ( .D(g25627), .SI(g3961), .SE(test_se), .CLK(CK), .Q(
        g962), .QN(n5630) );
  SDFFX1 DFF_417_Q_reg ( .D(g34657), .SI(g962), .SE(test_se), .CLK(CK), .Q(
        g101), .QN() );
  SDFFX1 DFF_418_Q_reg ( .D(g8870), .SI(g101), .SE(test_se), .CLK(CK), .Q(
        g8918), .QN(DFF_418_n1) );
  SDFFX1 DFF_419_Q_reg ( .D(g30552), .SI(g8918), .SE(test_se), .CLK(CK), .Q(
        g6625), .QN() );
  SDFFX1 DFF_420_Q_reg ( .D(g34979), .SI(g6625), .SE(test_se), .CLK(CK), .Q(
        n9332), .QN(DFF_420_n1) );
  SDFFX1 DFF_421_Q_reg ( .D(g30337), .SI(n9332), .SE(test_se), .CLK(CK), .Q(
        g1018), .QN() );
  SDFFX1 DFF_422_Q_reg ( .D(g24254), .SI(g1018), .SE(test_se), .CLK(CK), .Q(
        g17320), .QN() );
  SDFFX1 DFF_423_Q_reg ( .D(g24277), .SI(g17320), .SE(test_se), .CLK(CK), .Q(
        g4045), .QN() );
  SDFFX1 DFF_424_Q_reg ( .D(g29237), .SI(g4045), .SE(test_se), .CLK(CK), .Q(
        g1467), .QN(n5693) );
  SDFFX1 DFF_425_Q_reg ( .D(g30378), .SI(g1467), .SE(test_se), .CLK(CK), .Q(
        g2461), .QN(n5840) );
  SDFFX1 DFF_428_Q_reg ( .D(g33019), .SI(g2461), .SE(test_se), .CLK(CK), .Q(
        test_so30), .QN(n5300) );
  SDFFX1 DFF_429_Q_reg ( .D(g33623), .SI(test_si31), .SE(test_se), .CLK(CK), 
        .Q(g5990), .QN(n5589) );
  SDFFX1 DFF_431_Q_reg ( .D(g29235), .SI(g5990), .SE(test_se), .CLK(CK), .Q(
        g1256), .QN(n5558) );
  SDFFX1 DFF_432_Q_reg ( .D(g31902), .SI(g1256), .SE(test_se), .CLK(CK), .Q(
        g5029), .QN(n5601) );
  SDFFX1 DFF_433_Q_reg ( .D(g29306), .SI(g5029), .SE(test_se), .CLK(CK), .Q(
        g6519), .QN(n5806) );
  SDFFX1 DFF_434_Q_reg ( .D(g25689), .SI(g6519), .SE(test_se), .CLK(CK), .Q(
        g4169), .QN(n5729) );
  SDFFX1 DFF_435_Q_reg ( .D(g33978), .SI(g4169), .SE(test_se), .CLK(CK), .Q(
        g1816), .QN() );
  SDFFX1 DFF_436_Q_reg ( .D(g26970), .SI(g1816), .SE(test_se), .CLK(CK), .Q(
        g4369), .QN() );
  SDFFX1 DFF_439_Q_reg ( .D(g29278), .SI(g4369), .SE(test_se), .CLK(CK), .Q(
        g4578), .QN() );
  SDFFX1 DFF_440_Q_reg ( .D(g34253), .SI(g4578), .SE(test_se), .CLK(CK), .Q(
        g4459), .QN(n5765) );
  SDFFX1 DFF_441_Q_reg ( .D(g29272), .SI(g4459), .SE(test_se), .CLK(CK), .Q(
        g3831), .QN(n5872) );
  SDFFX1 DFF_442_Q_reg ( .D(g33595), .SI(g3831), .SE(test_se), .CLK(CK), .Q(
        g2514), .QN() );
  SDFFX1 DFF_443_Q_reg ( .D(g33610), .SI(g2514), .SE(test_se), .CLK(CK), .Q(
        g3288), .QN(n5400) );
  SDFFX1 DFF_444_Q_reg ( .D(g33589), .SI(g3288), .SE(test_se), .CLK(CK), .Q(
        test_so31), .QN(n5279) );
  SDFFX1 DFF_445_Q_reg ( .D(g34605), .SI(test_si32), .SE(test_se), .CLK(CK), 
        .Q(g2145), .QN(n5307) );
  SDFFX1 DFF_446_Q_reg ( .D(g30350), .SI(g2145), .SE(test_se), .CLK(CK), .Q(
        g1700), .QN(n5417) );
  SDFFX1 DFF_447_Q_reg ( .D(g25611), .SI(g1700), .SE(test_se), .CLK(CK), .Q(
        g513), .QN(n5548) );
  SDFFX1 DFF_448_Q_reg ( .D(test_so9), .SI(g513), .SE(test_se), .CLK(CK), .Q(
        g2841), .QN(n5963) );
  SDFFX1 DFF_449_Q_reg ( .D(g33619), .SI(g2841), .SE(test_se), .CLK(CK), .Q(
        g5297), .QN(n5588) );
  SDFFX1 DFF_451_Q_reg ( .D(g34022), .SI(g5297), .SE(test_se), .CLK(CK), .Q(
        g2763), .QN() );
  SDFFX1 DFF_452_Q_reg ( .D(g34033), .SI(g2763), .SE(test_se), .CLK(CK), .Q(
        g4793), .QN(n5368) );
  SDFFX1 DFF_453_Q_reg ( .D(g34726), .SI(g4793), .SE(test_se), .CLK(CK), .Q(
        g952), .QN() );
  SDFFX1 DFF_454_Q_reg ( .D(g31870), .SI(g952), .SE(test_se), .CLK(CK), .Q(
        g1263), .QN(n5674) );
  SDFFX1 DFF_455_Q_reg ( .D(g33985), .SI(g1263), .SE(test_se), .CLK(CK), .Q(
        g1950), .QN() );
  SDFFX1 DFF_456_Q_reg ( .D(g29283), .SI(g1950), .SE(test_se), .CLK(CK), .Q(
        g5138), .QN(n5871) );
  SDFFX1 DFF_457_Q_reg ( .D(g34003), .SI(g5138), .SE(test_se), .CLK(CK), .Q(
        g2307), .QN(n5859) );
  SDFFX1 DFF_458_Q_reg ( .D(g9497), .SI(g2307), .SE(test_se), .CLK(CK), .Q(
        test_so32), .QN() );
  SDFFX1 DFF_460_Q_reg ( .D(g25677), .SI(test_si33), .SE(test_se), .CLK(CK), 
        .Q(g8398), .QN() );
  SDFFX1 DFF_461_Q_reg ( .D(g34463), .SI(g8398), .SE(test_se), .CLK(CK), .Q(
        g4664), .QN() );
  SDFFX1 DFF_462_Q_reg ( .D(g33006), .SI(g4664), .SE(test_se), .CLK(CK), .Q(
        g2223), .QN(n5406) );
  SDFFX1 DFF_463_Q_reg ( .D(g29292), .SI(g2223), .SE(test_se), .CLK(CK), .Q(
        g5808), .QN(n5749) );
  SDFFX1 DFF_464_Q_reg ( .D(g30557), .SI(g5808), .SE(test_se), .CLK(CK), .Q(
        g6645), .QN() );
  SDFFX1 DFF_465_Q_reg ( .D(g33989), .SI(g6645), .SE(test_se), .CLK(CK), .Q(
        g2016), .QN(n5852) );
  SDFFX1 DFF_467_Q_reg ( .D(g33033), .SI(g2016), .SE(test_se), .CLK(CK), .Q(
        g3873), .QN(n5387) );
  SDFFX1 DFF_468_Q_reg ( .D(g11388), .SI(g3873), .SE(test_se), .CLK(CK), .Q(
        g13926), .QN(n5699) );
  SDFFX1 DFF_469_Q_reg ( .D(g34005), .SI(g13926), .SE(test_se), .CLK(CK), .Q(
        g2315), .QN(n5802) );
  SDFFX1 DFF_470_Q_reg ( .D(g26932), .SI(g2315), .SE(test_se), .CLK(CK), .Q(
        g2811), .QN() );
  SDFFX1 DFF_471_Q_reg ( .D(g30516), .SI(g2811), .SE(test_se), .CLK(CK), .Q(
        g5957), .QN() );
  SDFFX1 DFF_472_Q_reg ( .D(g33575), .SI(g5957), .SE(test_se), .CLK(CK), .Q(
        g2047), .QN(n5831) );
  SDFFX1 DFF_473_Q_reg ( .D(g33032), .SI(g2047), .SE(test_se), .CLK(CK), .Q(
        test_so33), .QN(n5648) );
  SDFFX1 DFF_474_Q_reg ( .D(g14779), .SI(test_si34), .SE(test_se), .CLK(CK), 
        .Q(g17760), .QN() );
  SDFFX1 DFF_476_Q_reg ( .D(g30486), .SI(g17760), .SE(test_se), .CLK(CK), .Q(
        g5575), .QN() );
  SDFFX1 DFF_477_Q_reg ( .D(g34974), .SI(g5575), .SE(test_se), .CLK(CK), .Q(
        n9327), .QN(DFF_477_n1) );
  SDFFX1 DFF_478_Q_reg ( .D(g25678), .SI(n9327), .SE(test_se), .CLK(CK), .Q(
        g3752), .QN(n5994) );
  SDFFX1 DFF_479_Q_reg ( .D(g30440), .SI(g3752), .SE(test_se), .CLK(CK), .Q(
        g3917), .QN() );
  SDFFX1 DFF_480_Q_reg ( .D(g11447), .SI(g3917), .SE(test_se), .CLK(CK), .Q(
        g8783), .QN(DFF_480_n1) );
  SDFFX1 DFF_481_Q_reg ( .D(g12923), .SI(g8783), .SE(test_se), .CLK(CK), .Q(
        g1585), .QN(n5757) );
  SDFFX1 DFF_482_Q_reg ( .D(g26949), .SI(g1585), .SE(test_se), .CLK(CK), .Q(
        g4388), .QN() );
  SDFFX1 DFF_483_Q_reg ( .D(g30530), .SI(g4388), .SE(test_se), .CLK(CK), .Q(
        g6275), .QN() );
  SDFFX1 DFF_484_Q_reg ( .D(g30542), .SI(g6275), .SE(test_se), .CLK(CK), .Q(
        g6311), .QN() );
  SDFFX1 DFF_485_Q_reg ( .D(g8915), .SI(g6311), .SE(test_se), .CLK(CK), .Q(
        g8916), .QN() );
  SDFFX1 DFF_486_Q_reg ( .D(g25624), .SI(g8916), .SE(test_se), .CLK(CK), .Q(
        g1041), .QN() );
  SDFFX1 DFF_487_Q_reg ( .D(g30383), .SI(g1041), .SE(test_se), .CLK(CK), .Q(
        test_so34), .QN(n5835) );
  SDFFX1 DFF_488_Q_reg ( .D(g33597), .SI(test_si35), .SE(test_se), .CLK(CK), 
        .Q(g2537), .QN(n5411) );
  SDFFX1 DFF_489_Q_reg ( .D(g34598), .SI(g2537), .SE(test_se), .CLK(CK), .Q(
        g21292), .QN(g30329) );
  SDFFX1 DFF_490_Q_reg ( .D(g26957), .SI(g21292), .SE(test_se), .CLK(CK), .Q(
        g4430), .QN() );
  SDFFX1 DFF_491_Q_reg ( .D(g26967), .SI(g4430), .SE(test_se), .CLK(CK), .Q(
        n9325), .QN(DFF_491_n1) );
  SDFFX1 DFF_493_Q_reg ( .D(g28102), .SI(n9325), .SE(test_se), .CLK(CK), .Q(
        g4826), .QN() );
  SDFFX1 DFF_494_Q_reg ( .D(g30524), .SI(g4826), .SE(test_se), .CLK(CK), .Q(
        g6239), .QN() );
  SDFFX1 DFF_496_Q_reg ( .D(g26903), .SI(g6239), .SE(test_se), .CLK(CK), .Q(
        g232), .QN() );
  SDFFX1 DFF_497_Q_reg ( .D(g30475), .SI(g232), .SE(test_se), .CLK(CK), .Q(
        g5268), .QN() );
  SDFFX1 DFF_498_Q_reg ( .D(g34647), .SI(g5268), .SE(test_se), .CLK(CK), .Q(
        g6545), .QN(n5497) );
  SDFFX1 DFF_499_Q_reg ( .D(g30377), .SI(g6545), .SE(test_se), .CLK(CK), .Q(
        n9324), .QN(n5314) );
  SDFFX1 DFF_500_Q_reg ( .D(g33553), .SI(n9324), .SE(test_se), .CLK(CK), .Q(
        g1772), .QN(n5504) );
  SDFFX1 DFF_502_Q_reg ( .D(g31903), .SI(g1772), .SE(test_se), .CLK(CK), .Q(
        g5052), .QN(n5607) );
  SDFFX1 DFF_503_Q_reg ( .D(g25715), .SI(g5052), .SE(test_se), .CLK(CK), .Q(
        g9615), .QN() );
  SDFFX1 DFF_504_Q_reg ( .D(g33984), .SI(test_si36), .SE(test_se), .CLK(CK), 
        .Q(g1890), .QN(n5799) );
  SDFFX1 DFF_505_Q_reg ( .D(g33602), .SI(g1890), .SE(test_se), .CLK(CK), .Q(
        g2629), .QN(n5521) );
  SDFFX1 DFF_506_Q_reg ( .D(g28045), .SI(g2629), .SE(test_se), .CLK(CK), .Q(
        g572), .QN(n5337) );
  SDFFX1 DFF_507_Q_reg ( .D(g34603), .SI(g572), .SE(test_se), .CLK(CK), .Q(
        g2130), .QN(n5487) );
  SDFFX1 DFF_508_Q_reg ( .D(g33035), .SI(g2130), .SE(test_se), .CLK(CK), .Q(
        g4108), .QN(n5715) );
  SDFFX1 DFF_509_Q_reg ( .D(g9251), .SI(g4108), .SE(test_se), .CLK(CK), .Q(
        g4308), .QN() );
  SDFFX1 DFF_510_Q_reg ( .D(g24208), .SI(g4308), .SE(test_se), .CLK(CK), .Q(
        g475), .QN() );
  SDFFX1 DFF_511_Q_reg ( .D(g8416), .SI(g475), .SE(test_se), .CLK(CK), .Q(g990), .QN(n5622) );
  SDFFX1 DFF_512_Q_reg ( .D(g34971), .SI(g990), .SE(test_se), .CLK(CK), .Q(g31), .QN(n5469) );
  SDFFX1 DFF_514_Q_reg ( .D(g34970), .SI(g31), .SE(test_se), .CLK(CK), .Q(
        n9322), .QN(DFF_514_n1) );
  SDFFX1 DFF_515_Q_reg ( .D(g24213), .SI(n9322), .SE(test_se), .CLK(CK), .Q(
        g12184), .QN() );
  SDFFX1 DFF_517_Q_reg ( .D(g33614), .SI(g12184), .SE(test_se), .CLK(CK), .Q(
        g3990), .QN(n5594) );
  SDFFX1 DFF_519_Q_reg ( .D(g33060), .SI(g3990), .SE(test_se), .CLK(CK), .Q(
        test_so36), .QN(n5565) );
  SDFFX1 DFF_520_Q_reg ( .D(g30362), .SI(test_si37), .SE(test_se), .CLK(CK), 
        .Q(g1992), .QN(n5890) );
  SDFFX1 DFF_522_Q_reg ( .D(g33023), .SI(g1992), .SE(test_se), .CLK(CK), .Q(
        g3171), .QN(n5603) );
  SDFFX1 DFF_524_Q_reg ( .D(g26898), .SI(g3171), .SE(test_se), .CLK(CK), .Q(
        g812), .QN(n5733) );
  SDFFX1 DFF_525_Q_reg ( .D(g25618), .SI(g812), .SE(test_se), .CLK(CK), .Q(
        g832), .QN() );
  SDFFX1 DFF_526_Q_reg ( .D(g30518), .SI(g832), .SE(test_se), .CLK(CK), .Q(
        g5897), .QN() );
  SDFFX1 DFF_527_Q_reg ( .D(g25688), .SI(g5897), .SE(test_se), .CLK(CK), .Q(
        g25689), .QN() );
  SDFFX1 DFF_528_Q_reg ( .D(g4570), .SI(g25689), .SE(test_se), .CLK(CK), .Q(
        g4571), .QN() );
  SDFFX1 DFF_529_Q_reg ( .D(g11349), .SI(g4571), .SE(test_se), .CLK(CK), .Q(
        g13895), .QN(n5702) );
  SDFFX1 DFF_530_Q_reg ( .D(g26959), .SI(g13895), .SE(test_se), .CLK(CK), .Q(
        g4455), .QN() );
  SDFFX1 DFF_531_Q_reg ( .D(g34801), .SI(g4455), .SE(test_se), .CLK(CK), .Q(
        g2902), .QN() );
  SDFFX1 DFF_532_Q_reg ( .D(g26884), .SI(g2902), .SE(test_se), .CLK(CK), .Q(
        g333), .QN() );
  SDFFX1 DFF_533_Q_reg ( .D(g25600), .SI(g333), .SE(test_se), .CLK(CK), .Q(
        g168), .QN(n5606) );
  SDFFX1 DFF_534_Q_reg ( .D(g26933), .SI(g168), .SE(test_se), .CLK(CK), .Q(
        test_so37), .QN() );
  SDFFX1 DFF_535_Q_reg ( .D(g28066), .SI(test_si38), .SE(test_se), .CLK(CK), 
        .Q(g3684), .QN(n5881) );
  SDFFX1 DFF_536_Q_reg ( .D(g33612), .SI(g3684), .SE(test_se), .CLK(CK), .Q(
        g3639), .QN(n5591) );
  SDFFX1 DFF_537_Q_reg ( .D(g17787), .SI(g3639), .SE(test_se), .CLK(CK), .Q(
        g14597), .QN(n5579) );
  SDFFX1 DFF_538_Q_reg ( .D(g24268), .SI(g14597), .SE(test_se), .CLK(CK), .Q(
        g3338), .QN(n5527) );
  SDFFX1 DFF_539_Q_reg ( .D(g25716), .SI(g3338), .SE(test_se), .CLK(CK), .Q(
        g5406), .QN(n5992) );
  SDFFX1 DFF_541_Q_reg ( .D(g26906), .SI(g5406), .SE(test_se), .CLK(CK), .Q(
        g269), .QN() );
  SDFFX1 DFF_542_Q_reg ( .D(g24203), .SI(g269), .SE(test_se), .CLK(CK), .Q(
        g401), .QN() );
  SDFFX1 DFF_543_Q_reg ( .D(g24346), .SI(g401), .SE(test_se), .CLK(CK), .Q(
        g6040), .QN() );
  SDFFX1 DFF_544_Q_reg ( .D(g24207), .SI(g6040), .SE(test_se), .CLK(CK), .Q(
        g441), .QN() );
  SDFFX1 DFF_545_Q_reg ( .D(g25701), .SI(g441), .SE(test_se), .CLK(CK), .Q(
        g9553), .QN(n5690) );
  SDFFX1 DFF_546_Q_reg ( .D(g29269), .SI(g9553), .SE(test_se), .CLK(CK), .Q(
        g3808), .QN(n5745) );
  SDFFX1 DFF_547_Q_reg ( .D(g34976), .SI(g3808), .SE(test_se), .CLK(CK), .Q(g9), .QN(n5468) );
  SDFFX1 DFF_549_Q_reg ( .D(g34255), .SI(g9), .SE(test_se), .CLK(CK), .Q(
        test_so38), .QN() );
  SDFFX1 DFF_550_Q_reg ( .D(g30450), .SI(test_si39), .SE(test_se), .CLK(CK), 
        .Q(g3957), .QN() );
  SDFFX1 DFF_551_Q_reg ( .D(g30456), .SI(g3957), .SE(test_se), .CLK(CK), .Q(
        g4093), .QN(n5340) );
  SDFFX1 DFF_552_Q_reg ( .D(g32991), .SI(g4093), .SE(test_se), .CLK(CK), .Q(
        g1760), .QN(n5602) );
  SDFFX1 DFF_554_Q_reg ( .D(g24348), .SI(g1760), .SE(test_se), .CLK(CK), .Q(
        g12422), .QN(n5437) );
  SDFFX1 DFF_555_Q_reg ( .D(g34249), .SI(g12422), .SE(test_se), .CLK(CK), .Q(
        g160), .QN(n5843) );
  SDFFX1 DFF_558_Q_reg ( .D(g30371), .SI(g160), .SE(test_se), .CLK(CK), .Q(
        g2279), .QN(n5778) );
  SDFFX1 DFF_559_Q_reg ( .D(g29268), .SI(g2279), .SE(test_se), .CLK(CK), .Q(
        g3498), .QN(n5740) );
  SDFFX1 DFF_560_Q_reg ( .D(g29224), .SI(g3498), .SE(test_se), .CLK(CK), .Q(
        g586), .QN(n5336) );
  SDFFX1 DFF_561_Q_reg ( .D(g14189), .SI(g586), .SE(test_se), .CLK(CK), .Q(
        g14201), .QN() );
  SDFFX1 DFF_562_Q_reg ( .D(g33017), .SI(g14201), .SE(test_se), .CLK(CK), .Q(
        g2619), .QN(n5508) );
  SDFFX1 DFF_563_Q_reg ( .D(g30339), .SI(g2619), .SE(test_se), .CLK(CK), .Q(
        g1183), .QN(n5599) );
  SDFFX1 DFF_564_Q_reg ( .D(g33967), .SI(g1183), .SE(test_se), .CLK(CK), .Q(
        g1608), .QN(n5792) );
  SDFFX1 DFF_565_Q_reg ( .D(g8784), .SI(g1608), .SE(test_se), .CLK(CK), .Q(
        g8785), .QN() );
  SDFFX1 DFF_566_Q_reg ( .D(g17519), .SI(test_si40), .SE(test_se), .CLK(CK), 
        .Q(g17577), .QN() );
  SDFFX1 DFF_567_Q_reg ( .D(g33559), .SI(g17577), .SE(test_se), .CLK(CK), .Q(
        g1779), .QN(n5830) );
  SDFFX1 DFF_568_Q_reg ( .D(g29255), .SI(g1779), .SE(test_se), .CLK(CK), .Q(
        g2652), .QN() );
  SDFFX1 DFF_570_Q_reg ( .D(g30368), .SI(g2652), .SE(test_se), .CLK(CK), .Q(
        g2193), .QN(n5839) );
  SDFFX1 DFF_571_Q_reg ( .D(g30375), .SI(g2193), .SE(test_se), .CLK(CK), .Q(
        g2393), .QN(n5421) );
  SDFFX1 DFF_573_Q_reg ( .D(g28052), .SI(g2393), .SE(test_se), .CLK(CK), .Q(
        g661), .QN() );
  SDFFX1 DFF_574_Q_reg ( .D(g28089), .SI(g661), .SE(test_se), .CLK(CK), .Q(
        g4950), .QN(n5772) );
  SDFFX1 DFF_575_Q_reg ( .D(g33055), .SI(g4950), .SE(test_se), .CLK(CK), .Q(
        g5535), .QN(n5566) );
  SDFFX1 DFF_576_Q_reg ( .D(g30392), .SI(g5535), .SE(test_se), .CLK(CK), .Q(
        g2834), .QN(g30330) );
  SDFFX1 DFF_577_Q_reg ( .D(g30343), .SI(g2834), .SE(test_se), .CLK(CK), .Q(
        g1361), .QN() );
  SDFFX1 DFF_579_Q_reg ( .D(g30523), .SI(g1361), .SE(test_se), .CLK(CK), .Q(
        g6235), .QN() );
  SDFFX1 DFF_580_Q_reg ( .D(g24233), .SI(g6235), .SE(test_se), .CLK(CK), .Q(
        g1146), .QN(n5851) );
  SDFFX1 DFF_581_Q_reg ( .D(g33018), .SI(g1146), .SE(test_se), .CLK(CK), .Q(
        test_so40), .QN(n5277) );
  SDFFX1 DFF_582_Q_reg ( .D(g32976), .SI(test_si41), .SE(test_se), .CLK(CK), 
        .Q(g150), .QN(n5676) );
  SDFFX1 DFF_583_Q_reg ( .D(g30349), .SI(g150), .SE(test_se), .CLK(CK), .Q(
        g1696), .QN(n5628) );
  SDFFX1 DFF_584_Q_reg ( .D(g33067), .SI(g1696), .SE(test_se), .CLK(CK), .Q(
        g6555), .QN() );
  SDFFX1 DFF_585_Q_reg ( .D(g26900), .SI(g6555), .SE(test_se), .CLK(CK), .Q(
        g14189), .QN() );
  SDFFX1 DFF_587_Q_reg ( .D(g33034), .SI(g14189), .SE(test_se), .CLK(CK), .Q(
        g3881), .QN(n5564) );
  SDFFX1 DFF_588_Q_reg ( .D(g30551), .SI(g3881), .SE(test_se), .CLK(CK), .Q(
        g6621), .QN() );
  SDFFX1 DFF_589_Q_reg ( .D(g25667), .SI(g6621), .SE(test_se), .CLK(CK), .Q(
        g3470), .QN(n5424) );
  SDFFX1 DFF_590_Q_reg ( .D(g30452), .SI(g3470), .SE(test_se), .CLK(CK), .Q(
        g3897), .QN() );
  SDFFX1 DFF_593_Q_reg ( .D(g34719), .SI(g518), .SE(test_se), .CLK(CK), .Q(
        g538), .QN(n5491) );
  SDFFX1 DFF_594_Q_reg ( .D(g33607), .SI(g538), .SE(test_se), .CLK(CK), .Q(
        g2606), .QN(n5311) );
  SDFFX1 DFF_595_Q_reg ( .D(g26923), .SI(g2606), .SE(test_se), .CLK(CK), .Q(
        g1472), .QN(n5290) );
  SDFFX1 DFF_597_Q_reg ( .D(g24211), .SI(g1472), .SE(test_se), .CLK(CK), .Q(
        test_so41), .QN(n5486) );
  SDFFX1 DFF_598_Q_reg ( .D(g33050), .SI(test_si42), .SE(test_se), .CLK(CK), 
        .Q(g5188), .QN(n5567) );
  SDFFX1 DFF_599_Q_reg ( .D(g24341), .SI(g5188), .SE(test_se), .CLK(CK), .Q(
        g5689), .QN(n5529) );
  SDFFX1 DFF_600_Q_reg ( .D(g19334), .SI(g5689), .SE(test_se), .CLK(CK), .Q(
        g13259), .QN() );
  SDFFX1 DFF_601_Q_reg ( .D(g24201), .SI(g13259), .SE(test_se), .CLK(CK), .Q(
        g405), .QN() );
  SDFFX1 DFF_602_Q_reg ( .D(g30463), .SI(g405), .SE(test_se), .CLK(CK), .Q(
        g5216), .QN() );
  SDFFX1 DFF_603_Q_reg ( .D(g9743), .SI(g5216), .SE(test_se), .CLK(CK), .Q(
        g6494), .QN() );
  SDFFX1 DFF_604_Q_reg ( .D(g34464), .SI(g6494), .SE(test_se), .CLK(CK), .Q(
        g4669), .QN() );
  SDFFX1 DFF_606_Q_reg ( .D(g24243), .SI(g4669), .SE(test_se), .CLK(CK), .Q(
        g996), .QN() );
  SDFFX1 DFF_607_Q_reg ( .D(g24335), .SI(g996), .SE(test_se), .CLK(CK), .Q(
        g4531), .QN() );
  SDFFX1 DFF_608_Q_reg ( .D(g34611), .SI(g4531), .SE(test_se), .CLK(CK), .Q(
        g2860), .QN() );
  SDFFX1 DFF_609_Q_reg ( .D(g34262), .SI(g2860), .SE(test_se), .CLK(CK), .Q(
        g4743), .QN(n5876) );
  SDFFX1 DFF_610_Q_reg ( .D(g30546), .SI(g4743), .SE(test_se), .CLK(CK), .Q(
        g6593), .QN() );
  SDFFX1 DFF_612_Q_reg ( .D(g25591), .SI(g6593), .SE(test_se), .CLK(CK), .Q(
        g8291), .QN() );
  SDFFX1 DFF_613_Q_reg ( .D(g7257), .SI(test_si43), .SE(test_se), .CLK(CK), 
        .Q(g4411), .QN() );
  SDFFX1 DFF_614_Q_reg ( .D(g30347), .SI(g4411), .SE(test_se), .CLK(CK), .Q(
        g1413), .QN() );
  SDFFX1 DFF_615_Q_reg ( .D(test_so38), .SI(g1413), .SE(test_se), .CLK(CK), 
        .Q(g26960), .QN() );
  SDFFX1 DFF_616_Q_reg ( .D(g17577), .SI(g26960), .SE(test_se), .CLK(CK), .Q(
        g13039), .QN() );
  SDFFX1 DFF_617_Q_reg ( .D(g30556), .SI(g13039), .SE(test_se), .CLK(CK), .Q(
        g6641), .QN() );
  SDFFX1 DFF_619_Q_reg ( .D(g34970), .SI(g6641), .SE(test_se), .CLK(CK), .Q(g6), .QN() );
  SDFFX1 DFF_620_Q_reg ( .D(g33562), .SI(g6), .SE(test_se), .CLK(CK), .Q(g1936), .QN(n5534) );
  SDFFX1 DFF_621_Q_reg ( .D(n1278), .SI(g1936), .SE(test_se), .CLK(CK), .Q(g55), .QN() );
  SDFFX1 DFF_622_Q_reg ( .D(g25610), .SI(g55), .SE(test_se), .CLK(CK), .Q(g504), .QN(n5519) );
  SDFFX1 DFF_623_Q_reg ( .D(g33015), .SI(g504), .SE(test_se), .CLK(CK), .Q(
        g2587), .QN(n5372) );
  SDFFX1 DFF_624_Q_reg ( .D(g31896), .SI(g2587), .SE(test_se), .CLK(CK), .Q(
        g4480), .QN() );
  SDFFX1 DFF_625_Q_reg ( .D(g34004), .SI(g4480), .SE(test_se), .CLK(CK), .Q(
        n9314), .QN(n5687) );
  SDFFX1 DFF_626_Q_reg ( .D(g30428), .SI(n9314), .SE(test_se), .CLK(CK), .Q(
        test_so43), .QN() );
  SDFFX1 DFF_627_Q_reg ( .D(g30485), .SI(test_si44), .SE(test_se), .CLK(CK), 
        .Q(g5571), .QN() );
  SDFFX1 DFF_628_Q_reg ( .D(g30422), .SI(g5571), .SE(test_se), .CLK(CK), .Q(
        g3578), .QN() );
  SDFFX1 DFF_630_Q_reg ( .D(g25714), .SI(g3578), .SE(test_se), .CLK(CK), .Q(
        g9555), .QN(n5720) );
  SDFFX1 DFF_632_Q_reg ( .D(g29294), .SI(g9555), .SE(test_se), .CLK(CK), .Q(
        g5827), .QN(n5809) );
  SDFFX1 DFF_633_Q_reg ( .D(g30423), .SI(g5827), .SE(test_se), .CLK(CK), .Q(
        g3582), .QN() );
  SDFFX1 DFF_634_Q_reg ( .D(g30529), .SI(g3582), .SE(test_se), .CLK(CK), .Q(
        g6271), .QN() );
  SDFFX1 DFF_635_Q_reg ( .D(g34028), .SI(g6271), .SE(test_se), .CLK(CK), .Q(
        g4688), .QN(n5656) );
  SDFFX1 DFF_637_Q_reg ( .D(g33587), .SI(g4688), .SE(test_se), .CLK(CK), .Q(
        g2380), .QN() );
  SDFFX1 DFF_638_Q_reg ( .D(g30460), .SI(g2380), .SE(test_se), .CLK(CK), .Q(
        g5196), .QN() );
  SDFFX1 DFF_640_Q_reg ( .D(g30401), .SI(g5196), .SE(test_se), .CLK(CK), .Q(
        g3227), .QN() );
  SDFFX1 DFF_641_Q_reg ( .D(g33990), .SI(g3227), .SE(test_se), .CLK(CK), .Q(
        n9312), .QN(n5683) );
  SDFFX1 DFF_642_Q_reg ( .D(g16693), .SI(n9312), .SE(test_se), .CLK(CK), .Q(
        g14518), .QN() );
  SDFFX1 DFF_643_Q_reg ( .D(g17291), .SI(g14518), .SE(test_se), .CLK(CK), .Q(
        g17316), .QN() );
  SDFFX1 DFF_644_Q_reg ( .D(g29309), .SI(test_si45), .SE(test_se), .CLK(CK), 
        .Q(g6541), .QN(n5739) );
  SDFFX1 DFF_645_Q_reg ( .D(g30411), .SI(g6541), .SE(test_se), .CLK(CK), .Q(
        g3203), .QN() );
  SDFFX1 DFF_646_Q_reg ( .D(g33546), .SI(g3203), .SE(test_se), .CLK(CK), .Q(
        g1668), .QN(n5598) );
  SDFFX1 DFF_647_Q_reg ( .D(g28085), .SI(g1668), .SE(test_se), .CLK(CK), .Q(
        g4760), .QN(n5775) );
  SDFFX1 DFF_648_Q_reg ( .D(g26904), .SI(g4760), .SE(test_se), .CLK(CK), .Q(
        g262), .QN() );
  SDFFX1 DFF_649_Q_reg ( .D(g33556), .SI(g262), .SE(test_se), .CLK(CK), .Q(
        g1840), .QN(n5451) );
  SDFFX1 DFF_651_Q_reg ( .D(g25722), .SI(g1840), .SE(test_se), .CLK(CK), .Q(
        g5467), .QN() );
  SDFFX1 DFF_652_Q_reg ( .D(g25605), .SI(g5467), .SE(test_se), .CLK(CK), .Q(
        g460), .QN() );
  SDFFX1 DFF_653_Q_reg ( .D(g33062), .SI(g460), .SE(test_se), .CLK(CK), .Q(
        g6209), .QN() );
  SDFFX1 DFF_654_Q_reg ( .D(g26893), .SI(g6209), .SE(test_se), .CLK(CK), .Q(
        g20763), .QN() );
  SDFFX1 DFF_655_Q_reg ( .D(g12238), .SI(g20763), .SE(test_se), .CLK(CK), .Q(
        g14662), .QN(n5704) );
  SDFFX1 DFF_656_Q_reg ( .D(g28050), .SI(g14662), .SE(test_se), .CLK(CK), .Q(
        g655), .QN() );
  SDFFX1 DFF_657_Q_reg ( .D(g34626), .SI(g655), .SE(test_se), .CLK(CK), .Q(
        test_so45), .QN(n5496) );
  SDFFX1 DFF_658_Q_reg ( .D(g33583), .SI(test_si46), .SE(test_se), .CLK(CK), 
        .Q(g2204), .QN(n5620) );
  SDFFX1 DFF_659_Q_reg ( .D(g30472), .SI(g2204), .SE(test_se), .CLK(CK), .Q(
        g5256), .QN() );
  SDFFX1 DFF_660_Q_reg ( .D(g34454), .SI(g5256), .SE(test_se), .CLK(CK), .Q(
        g4608), .QN(n5274) );
  SDFFX1 DFF_661_Q_reg ( .D(g34850), .SI(g4608), .SE(test_se), .CLK(CK), .Q(
        g794), .QN(n5291) );
  SDFFX1 DFF_662_Q_reg ( .D(g16955), .SI(g794), .SE(test_se), .CLK(CK), .Q(
        g13906), .QN(n5583) );
  SDFFX1 DFF_663_Q_reg ( .D(g10306), .SI(g13906), .SE(test_se), .CLK(CK), .Q(
        g4423), .QN() );
  SDFFX1 DFF_664_Q_reg ( .D(g24272), .SI(g4423), .SE(test_se), .CLK(CK), .Q(
        g3689), .QN(n5532) );
  SDFFX1 DFF_666_Q_reg ( .D(g17678), .SI(g3689), .SE(test_se), .CLK(CK), .Q(
        g5685), .QN() );
  SDFFX1 DFF_667_Q_reg ( .D(g24214), .SI(g5685), .SE(test_se), .CLK(CK), .Q(
        g703), .QN(n5821) );
  SDFFX1 DFF_669_Q_reg ( .D(g26909), .SI(g703), .SE(test_se), .CLK(CK), .Q(
        g862), .QN(n5682) );
  SDFFX1 DFF_670_Q_reg ( .D(g30406), .SI(g862), .SE(test_se), .CLK(CK), .Q(
        g3247), .QN() );
  SDFFX1 DFF_671_Q_reg ( .D(g33569), .SI(g3247), .SE(test_se), .CLK(CK), .Q(
        g2040), .QN(n5505) );
  SDFFX1 DFF_672_Q_reg ( .D(g25694), .SI(g2040), .SE(test_se), .CLK(CK), .Q(
        g8178), .QN(DFF_672_n1) );
  SDFFX1 DFF_673_Q_reg ( .D(g34628), .SI(test_si47), .SE(test_se), .CLK(CK), 
        .Q(g4146), .QN(n5981) );
  SDFFX1 DFF_674_Q_reg ( .D(g34458), .SI(g4146), .SE(test_se), .CLK(CK), .Q(
        g4633), .QN(n5844) );
  SDFFX1 DFF_675_Q_reg ( .D(g24240), .SI(g4633), .SE(test_se), .CLK(CK), .Q(
        g1157), .QN(n5304) );
  SDFFX1 DFF_677_Q_reg ( .D(g34634), .SI(g1157), .SE(test_se), .CLK(CK), .Q(
        g4732), .QN(n5296) );
  SDFFX1 DFF_678_Q_reg ( .D(g25700), .SI(g4732), .SE(test_se), .CLK(CK), .Q(
        g9497), .QN(n5689) );
  SDFFX1 DFF_679_Q_reg ( .D(g29293), .SI(g9497), .SE(test_se), .CLK(CK), .Q(
        g5817), .QN() );
  SDFFX1 DFF_681_Q_reg ( .D(g33009), .SI(g5817), .SE(test_se), .CLK(CK), .Q(
        g2351), .QN(n5511) );
  SDFFX1 DFF_682_Q_reg ( .D(g33603), .SI(g2351), .SE(test_se), .CLK(CK), .Q(
        g2648), .QN() );
  SDFFX1 DFF_683_Q_reg ( .D(g24355), .SI(g2648), .SE(test_se), .CLK(CK), .Q(
        g6736), .QN() );
  SDFFX1 DFF_684_Q_reg ( .D(g34268), .SI(g6736), .SE(test_se), .CLK(CK), .Q(
        g4944), .QN(n5875) );
  SDFFX1 DFF_685_Q_reg ( .D(g25691), .SI(g4944), .SE(test_se), .CLK(CK), .Q(
        g4072), .QN() );
  SDFFX1 DFF_686_Q_reg ( .D(g26890), .SI(g4072), .SE(test_se), .CLK(CK), .Q(
        g7540), .QN() );
  SDFFX1 DFF_687_Q_reg ( .D(g7260), .SI(g7540), .SE(test_se), .CLK(CK), .Q(
        test_so47), .QN() );
  SDFFX1 DFF_688_Q_reg ( .D(g29264), .SI(test_si48), .SE(test_se), .CLK(CK), 
        .Q(g3466), .QN() );
  SDFFX1 DFF_689_Q_reg ( .D(g28072), .SI(g3466), .SE(test_se), .CLK(CK), .Q(
        g4116), .QN() );
  SDFFX1 DFF_690_Q_reg ( .D(g31900), .SI(g4116), .SE(test_se), .CLK(CK), .Q(
        g5041), .QN(n5605) );
  SDFFX1 DFF_692_Q_reg ( .D(g26956), .SI(g5041), .SE(test_se), .CLK(CK), .Q(
        g4434), .QN() );
  SDFFX1 DFF_693_Q_reg ( .D(g29271), .SI(g4434), .SE(test_se), .CLK(CK), .Q(
        g3827), .QN(n5808) );
  SDFFX1 DFF_694_Q_reg ( .D(g29304), .SI(g3827), .SE(test_se), .CLK(CK), .Q(
        g6500), .QN(n5748) );
  SDFFX1 DFF_695_Q_reg ( .D(g13049), .SI(g6500), .SE(test_se), .CLK(CK), .Q(
        g17813), .QN() );
  SDFFX1 DFF_696_Q_reg ( .D(g29261), .SI(g17813), .SE(test_se), .CLK(CK), .Q(
        g3133), .QN(n5661) );
  SDFFX1 DFF_697_Q_reg ( .D(g28063), .SI(g3133), .SE(test_se), .CLK(CK), .Q(
        g3333), .QN() );
  SDFFX1 DFF_698_Q_reg ( .D(g13259), .SI(g3333), .SE(test_se), .CLK(CK), .Q(
        g979), .QN(n5320) );
  SDFFX1 DFF_699_Q_reg ( .D(g34027), .SI(g979), .SE(test_se), .CLK(CK), .Q(
        g4681), .QN() );
  SDFFX1 DFF_700_Q_reg ( .D(g33961), .SI(g4681), .SE(test_se), .CLK(CK), .Q(
        g298), .QN(n5675) );
  SDFFX1 DFF_702_Q_reg ( .D(g33604), .SI(g298), .SE(test_se), .CLK(CK), .Q(
        test_so48), .QN(n5759) );
  SDFFX1 DFF_704_Q_reg ( .D(g8788), .SI(test_si49), .SE(test_se), .CLK(CK), 
        .Q(g8789), .QN() );
  SDFFX1 DFF_705_Q_reg ( .D(g32995), .SI(g8789), .SE(test_se), .CLK(CK), .Q(
        g1894), .QN(n5374) );
  SDFFX1 DFF_706_Q_reg ( .D(g34624), .SI(g1894), .SE(test_se), .CLK(CK), .Q(
        g2988), .QN() );
  SDFFX1 DFF_707_Q_reg ( .D(g30415), .SI(g2988), .SE(test_se), .CLK(CK), .Q(
        g3538), .QN() );
  SDFFX1 DFF_708_Q_reg ( .D(g33536), .SI(g3538), .SE(test_se), .CLK(CK), .Q(
        g301), .QN() );
  SDFFX1 DFF_709_Q_reg ( .D(g26888), .SI(g301), .SE(test_se), .CLK(CK), .Q(
        n9306), .QN(DFF_709_n1) );
  SDFFX1 DFF_710_Q_reg ( .D(g28055), .SI(n9306), .SE(test_se), .CLK(CK), .Q(
        g827), .QN(n5728) );
  SDFFX1 DFF_711_Q_reg ( .D(g24238), .SI(g827), .SE(test_se), .CLK(CK), .Q(
        g17291), .QN() );
  SDFFX1 DFF_713_Q_reg ( .D(g33600), .SI(g17291), .SE(test_se), .CLK(CK), .Q(
        g2555), .QN(n5351) );
  SDFFX1 DFF_714_Q_reg ( .D(g28105), .SI(g2555), .SE(test_se), .CLK(CK), .Q(
        g5011), .QN() );
  SDFFX1 DFF_715_Q_reg ( .D(g34721), .SI(g5011), .SE(test_se), .CLK(CK), .Q(
        g199), .QN() );
  SDFFX1 DFF_716_Q_reg ( .D(g29307), .SI(g199), .SE(test_se), .CLK(CK), .Q(
        g6523), .QN(n5870) );
  SDFFX1 DFF_717_Q_reg ( .D(g30345), .SI(g6523), .SE(test_se), .CLK(CK), .Q(
        test_so49), .QN(n5542) );
  SDFFX1 DFF_718_Q_reg ( .D(g34453), .SI(test_si50), .SE(test_se), .CLK(CK), 
        .Q(g4601), .QN(n5365) );
  SDFFX1 DFF_719_Q_reg ( .D(g32980), .SI(g4601), .SE(test_se), .CLK(CK), .Q(
        g854), .QN(n5754) );
  SDFFX1 DFF_720_Q_reg ( .D(g29238), .SI(g854), .SE(test_se), .CLK(CK), .Q(
        g1484), .QN(n5865) );
  SDFFX1 DFF_721_Q_reg ( .D(g34639), .SI(g1484), .SE(test_se), .CLK(CK), .Q(
        g4922), .QN(n5346) );
  SDFFX1 DFF_722_Q_reg ( .D(g25695), .SI(g4922), .SE(test_se), .CLK(CK), .Q(
        g5080), .QN(n5893) );
  SDFFX1 DFF_723_Q_reg ( .D(g33057), .SI(g5080), .SE(test_se), .CLK(CK), .Q(
        g5863), .QN() );
  SDFFX1 DFF_724_Q_reg ( .D(g26969), .SI(g5863), .SE(test_se), .CLK(CK), .Q(
        g4581), .QN(n5670) );
  SDFFX1 DFF_726_Q_reg ( .D(g29253), .SI(g4581), .SE(test_se), .CLK(CK), .Q(
        g2518), .QN() );
  SDFFX1 DFF_727_Q_reg ( .D(g34021), .SI(g2518), .SE(test_se), .CLK(CK), .Q(
        g2567), .QN() );
  SDFFX1 DFF_728_Q_reg ( .D(g26895), .SI(g2567), .SE(test_se), .CLK(CK), .Q(
        g568), .QN(n5335) );
  SDFFX1 DFF_729_Q_reg ( .D(g30413), .SI(g568), .SE(test_se), .CLK(CK), .Q(
        g3263), .QN() );
  SDFFX1 DFF_730_Q_reg ( .D(g30549), .SI(g3263), .SE(test_se), .CLK(CK), .Q(
        g6613), .QN() );
  SDFFX1 DFF_731_Q_reg ( .D(g24347), .SI(g6613), .SE(test_se), .CLK(CK), .Q(
        test_so50), .QN() );
  SDFFX1 DFF_732_Q_reg ( .D(g25758), .SI(test_si51), .SE(test_se), .CLK(CK), 
        .Q(g6444), .QN(n5990) );
  SDFFX1 DFF_733_Q_reg ( .D(g34808), .SI(g6444), .SE(test_se), .CLK(CK), .Q(
        g2965), .QN() );
  SDFFX1 DFF_734_Q_reg ( .D(g30501), .SI(g2965), .SE(test_se), .CLK(CK), .Q(
        g5857), .QN(n5573) );
  SDFFX1 DFF_735_Q_reg ( .D(g33969), .SI(g5857), .SE(test_se), .CLK(CK), .Q(
        n9303), .QN(n5587) );
  SDFFX1 DFF_736_Q_reg ( .D(g34440), .SI(n9303), .SE(test_se), .CLK(CK), .Q(
        g890), .QN(n5305) );
  SDFFX1 DFF_737_Q_reg ( .D(g17607), .SI(g890), .SE(test_se), .CLK(CK), .Q(
        g17646), .QN() );
  SDFFX1 DFF_738_Q_reg ( .D(g30433), .SI(g17646), .SE(test_se), .CLK(CK), .Q(
        g3562), .QN() );
  SDFFX1 DFF_739_Q_reg ( .D(g21900), .SI(g3562), .SE(test_se), .CLK(CK), .Q(
        g10122_Tj), .QN() );
  SDFFX1 DFF_740_Q_reg ( .D(g26921), .SI(g10122_Tj), .SE(test_se), .CLK(CK), .Q(
        g1404), .QN() );
  SDFFX1 DFF_742_Q_reg ( .D(g29270), .SI(g1404), .SE(test_se), .CLK(CK), .Q(
        g3817), .QN() );
  SDFFX1 DFF_743_Q_reg ( .D(n1485), .SI(g3817), .SE(test_se), .CLK(CK), .Q(
        n9302), .QN(n6010) );
  SDFFX1 DFF_744_Q_reg ( .D(g33038), .SI(n9302), .SE(test_se), .CLK(CK), .Q(
        g4501), .QN() );
  SDFFX1 DFF_745_Q_reg ( .D(g31865), .SI(g4501), .SE(test_se), .CLK(CK), .Q(
        test_so51), .QN() );
  SDFFX1 DFF_746_Q_reg ( .D(g26926), .SI(test_si52), .SE(test_se), .CLK(CK), 
        .Q(g2724), .QN(n5301) );
  SDFFX1 DFF_747_Q_reg ( .D(g28083), .SI(g2724), .SE(test_se), .CLK(CK), .Q(
        g4704), .QN(n5771) );
  SDFFX1 DFF_749_Q_reg ( .D(g34797), .SI(g22), .SE(test_se), .CLK(CK), .Q(
        g2878), .QN() );
  SDFFX1 DFF_750_Q_reg ( .D(g30478), .SI(g2878), .SE(test_se), .CLK(CK), .Q(
        g5220), .QN() );
  SDFFX1 DFF_751_Q_reg ( .D(g34724), .SI(g5220), .SE(test_se), .CLK(CK), .Q(
        g617), .QN(n5339) );
  SDFFX1 DFF_752_Q_reg ( .D(g24212), .SI(g617), .SE(test_se), .CLK(CK), .Q(
        g12368), .QN(n5485) );
  SDFFX1 DFF_753_Q_reg ( .D(g26883), .SI(g12368), .SE(test_se), .CLK(CK), .Q(
        g316), .QN() );
  SDFFX1 DFF_754_Q_reg ( .D(g32985), .SI(g316), .SE(test_se), .CLK(CK), .Q(
        g1277), .QN() );
  SDFFX1 DFF_755_Q_reg ( .D(g25761), .SI(g1277), .SE(test_se), .CLK(CK), .Q(
        g6513), .QN(n5426) );
  SDFFX1 DFF_756_Q_reg ( .D(g26886), .SI(g6513), .SE(test_se), .CLK(CK), .Q(
        g336), .QN(n5824) );
  SDFFX1 DFF_757_Q_reg ( .D(g34796), .SI(g336), .SE(test_se), .CLK(CK), .Q(
        g2882), .QN() );
  SDFFX1 DFF_758_Q_reg ( .D(g32982), .SI(g2882), .SE(test_se), .CLK(CK), .Q(
        test_so52), .QN() );
  SDFFX1 DFF_759_Q_reg ( .D(g33561), .SI(test_si53), .SE(test_se), .CLK(CK), 
        .Q(g1906), .QN(n5503) );
  SDFFX1 DFF_760_Q_reg ( .D(g26880), .SI(g1906), .SE(test_se), .CLK(CK), .Q(
        g305), .QN(n5282) );
  SDFFX1 DFF_761_Q_reg ( .D(g34975), .SI(g305), .SE(test_se), .CLK(CK), .Q(g8), 
        .QN() );
  SDFFX1 DFF_763_Q_reg ( .D(g26931), .SI(g8), .SE(test_se), .CLK(CK), .Q(g2799), .QN() );
  SDFFX1 DFF_764_Q_reg ( .D(g14147), .SI(g2799), .SE(test_se), .CLK(CK), .Q(
        g14167), .QN() );
  SDFFX1 DFF_765_Q_reg ( .D(g13039), .SI(g14167), .SE(test_se), .CLK(CK), .Q(
        g17787), .QN() );
  SDFFX1 DFF_766_Q_reg ( .D(g34641), .SI(g17787), .SE(test_se), .CLK(CK), .Q(
        g4912), .QN(n5297) );
  SDFFX1 DFF_767_Q_reg ( .D(g34629), .SI(g4912), .SE(test_se), .CLK(CK), .Q(
        g4157), .QN(n5983) );
  SDFFX1 DFF_768_Q_reg ( .D(g33598), .SI(g4157), .SE(test_se), .CLK(CK), .Q(
        g2541), .QN(n5461) );
  SDFFX1 DFF_769_Q_reg ( .D(g33576), .SI(g2541), .SE(test_se), .CLK(CK), .Q(
        g2153), .QN(n5356) );
  SDFFX1 DFF_770_Q_reg ( .D(g34720), .SI(g2153), .SE(test_se), .CLK(CK), .Q(
        g550), .QN() );
  SDFFX1 DFF_771_Q_reg ( .D(g26902), .SI(g550), .SE(test_se), .CLK(CK), .Q(
        g255), .QN() );
  SDFFX1 DFF_772_Q_reg ( .D(g29244), .SI(g255), .SE(test_se), .CLK(CK), .Q(
        test_so53), .QN() );
  SDFFX1 DFF_773_Q_reg ( .D(g30468), .SI(test_si54), .SE(test_se), .CLK(CK), 
        .Q(g5240), .QN() );
  SDFFX1 DFF_774_Q_reg ( .D(g26924), .SI(g5240), .SE(test_se), .CLK(CK), .Q(
        g1478), .QN(n5289) );
  SDFFX1 DFF_776_Q_reg ( .D(g33031), .SI(g1478), .SE(test_se), .CLK(CK), .Q(
        g3863), .QN() );
  SDFFX1 DFF_777_Q_reg ( .D(g29245), .SI(g3863), .SE(test_se), .CLK(CK), .Q(
        g1959), .QN() );
  SDFFX1 DFF_778_Q_reg ( .D(g29266), .SI(g1959), .SE(test_se), .CLK(CK), .Q(
        g3480), .QN(n5868) );
  SDFFX1 DFF_779_Q_reg ( .D(g30559), .SI(g3480), .SE(test_se), .CLK(CK), .Q(
        g6653), .QN() );
  SDFFX1 DFF_780_Q_reg ( .D(g14749), .SI(g6653), .SE(test_se), .CLK(CK), .Q(
        g17764), .QN() );
  SDFFX1 DFF_781_Q_reg ( .D(g34794), .SI(g17764), .SE(test_se), .CLK(CK), .Q(
        g2864), .QN(n5489) );
  SDFFX1 DFF_782_Q_reg ( .D(g28087), .SI(g2864), .SE(test_se), .CLK(CK), .Q(
        g4894), .QN(n5774) );
  SDFFX1 DFF_783_Q_reg ( .D(g14635), .SI(g4894), .SE(test_se), .CLK(CK), .Q(
        g17678), .QN() );
  SDFFX1 DFF_784_Q_reg ( .D(g30435), .SI(g17678), .SE(test_se), .CLK(CK), .Q(
        g3857), .QN(n5572) );
  SDFFX1 DFF_785_Q_reg ( .D(g16659), .SI(g3857), .SE(test_se), .CLK(CK), .Q(
        g16693), .QN() );
  SDFFX1 DFF_786_Q_reg ( .D(g25609), .SI(g16693), .SE(test_se), .CLK(CK), .Q(
        test_so54), .QN(n5481) );
  SDFFX1 DFF_788_Q_reg ( .D(g28057), .SI(test_si55), .SE(test_se), .CLK(CK), 
        .Q(g1002), .QN() );
  SDFFX1 DFF_789_Q_reg ( .D(g34439), .SI(g1002), .SE(test_se), .CLK(CK), .Q(
        g776), .QN(n5330) );
  SDFFX1 DFF_790_Q_reg ( .D(g34979), .SI(g776), .SE(test_se), .CLK(CK), .Q(g28), .QN(n5324) );
  SDFFX1 DFF_791_Q_reg ( .D(g10500), .SI(g28), .SE(test_se), .CLK(CK), .Q(
        g1236), .QN() );
  SDFFX1 DFF_792_Q_reg ( .D(g34260), .SI(g1236), .SE(test_se), .CLK(CK), .Q(
        g4646), .QN(n5712) );
  SDFFX1 DFF_793_Q_reg ( .D(g33012), .SI(g4646), .SE(test_se), .CLK(CK), .Q(
        g2476), .QN() );
  SDFFX1 DFF_794_Q_reg ( .D(g32989), .SI(g2476), .SE(test_se), .CLK(CK), .Q(
        g1657), .QN(n5525) );
  SDFFX1 DFF_795_Q_reg ( .D(g34006), .SI(g1657), .SE(test_se), .CLK(CK), .Q(
        g2375), .QN() );
  SDFFX1 DFF_796_Q_reg ( .D(g34783), .SI(g2375), .SE(test_se), .CLK(CK), .Q(
        g63), .QN() );
  SDFFX1 DFF_797_Q_reg ( .D(g14738), .SI(g63), .SE(test_se), .CLK(CK), .Q(
        g17739), .QN() );
  SDFFX1 DFF_798_Q_reg ( .D(g8719), .SI(g17739), .SE(test_se), .CLK(CK), .Q(
        g358), .QN() );
  SDFFX1 DFF_799_Q_reg ( .D(g26910), .SI(g358), .SE(test_se), .CLK(CK), .Q(
        g896), .QN(n5431) );
  SDFFX1 DFF_802_Q_reg ( .D(g28043), .SI(g896), .SE(test_se), .CLK(CK), .Q(
        test_so55), .QN(n5695) );
  SDFFX1 DFF_803_Q_reg ( .D(g33021), .SI(test_si56), .SE(test_se), .CLK(CK), 
        .Q(g3161), .QN() );
  SDFFX1 DFF_804_Q_reg ( .D(g29251), .SI(g3161), .SE(test_se), .CLK(CK), .Q(
        g2384), .QN() );
  SDFFX1 DFF_806_Q_reg ( .D(g12470), .SI(g2384), .SE(test_se), .CLK(CK), .Q(
        g14828), .QN(n5700) );
  SDFFX1 DFF_807_Q_reg ( .D(g34456), .SI(g14828), .SE(test_se), .CLK(CK), .Q(
        g4616), .QN(n5608) );
  SDFFX1 DFF_808_Q_reg ( .D(g26968), .SI(g4616), .SE(test_se), .CLK(CK), .Q(
        g4561), .QN() );
  SDFFX1 DFF_809_Q_reg ( .D(g33991), .SI(g4561), .SE(test_se), .CLK(CK), .Q(
        g2024), .QN(n5801) );
  SDFFX1 DFF_810_Q_reg ( .D(g8279), .SI(g2024), .SE(test_se), .CLK(CK), .Q(
        g3451), .QN() );
  SDFFX1 DFF_811_Q_reg ( .D(g26930), .SI(g3451), .SE(test_se), .CLK(CK), .Q(
        g2795), .QN() );
  SDFFX1 DFF_812_Q_reg ( .D(g34599), .SI(g2795), .SE(test_se), .CLK(CK), .Q(
        g613), .QN(n5474) );
  SDFFX1 DFF_813_Q_reg ( .D(g28082), .SI(g613), .SE(test_se), .CLK(CK), .Q(
        g4527), .QN() );
  SDFFX1 DFF_814_Q_reg ( .D(g33557), .SI(g4527), .SE(test_se), .CLK(CK), .Q(
        g1844), .QN(n5847) );
  SDFFX1 DFF_815_Q_reg ( .D(g30511), .SI(g1844), .SE(test_se), .CLK(CK), .Q(
        g5937), .QN() );
  SDFFX1 DFF_816_Q_reg ( .D(g33045), .SI(g5937), .SE(test_se), .CLK(CK), .Q(
        test_so56), .QN() );
  SDFFX1 DFF_818_Q_reg ( .D(g30379), .SI(test_si57), .SE(test_se), .CLK(CK), 
        .Q(g2523), .QN(n5281) );
  SDFFX1 DFF_819_Q_reg ( .D(g24267), .SI(g2523), .SE(test_se), .CLK(CK), .Q(
        g11349), .QN(n5436) );
  SDFFX1 DFF_820_Q_reg ( .D(g34020), .SI(g11349), .SE(test_se), .CLK(CK), .Q(
        g2643), .QN() );
  SDFFX1 DFF_822_Q_reg ( .D(g24249), .SI(g2643), .SE(test_se), .CLK(CK), .Q(
        g1489), .QN(n5850) );
  SDFFX1 DFF_824_Q_reg ( .D(g25592), .SI(g1489), .SE(test_se), .CLK(CK), .Q(
        g8358), .QN() );
  SDFFX1 DFF_825_Q_reg ( .D(g30382), .SI(g8358), .SE(test_se), .CLK(CK), .Q(
        n9295), .QN(n5625) );
  SDFFX1 DFF_826_Q_reg ( .D(g29285), .SI(n9295), .SE(test_se), .CLK(CK), .Q(
        g5156), .QN(n5734) );
  SDFFX1 DFF_828_Q_reg ( .D(g12919), .SI(g5156), .SE(test_se), .CLK(CK), .Q(
        g23683), .QN(n5526) );
  SDFFX1 DFF_829_Q_reg ( .D(g34975), .SI(g23683), .SE(test_se), .CLK(CK), .Q(
        n9294), .QN(DFF_829_n1) );
  SDFFX1 DFF_830_Q_reg ( .D(g25662), .SI(n9294), .SE(test_se), .CLK(CK), .Q(
        g8279), .QN(n5717) );
  SDFFX1 DFF_831_Q_reg ( .D(g21896), .SI(g8279), .SE(test_se), .CLK(CK), .Q(
        g8839), .QN() );
  SDFFX1 DFF_832_Q_reg ( .D(g33563), .SI(g8839), .SE(test_se), .CLK(CK), .Q(
        g1955), .QN() );
  SDFFX1 DFF_833_Q_reg ( .D(g33622), .SI(g1955), .SE(test_se), .CLK(CK), .Q(
        test_so57), .QN(n5394) );
  SDFFX1 DFF_835_Q_reg ( .D(g33582), .SI(test_si58), .SE(test_se), .CLK(CK), 
        .Q(g2273), .QN(n5458) );
  SDFFX1 DFF_836_Q_reg ( .D(g17871), .SI(g2273), .SE(test_se), .CLK(CK), .Q(
        g14749), .QN(n5584) );
  SDFFX1 DFF_837_Q_reg ( .D(g28086), .SI(g14749), .SE(test_se), .CLK(CK), .Q(
        g4771), .QN(n5769) );
  SDFFX1 DFF_838_Q_reg ( .D(g25744), .SI(g4771), .SE(test_se), .CLK(CK), .Q(
        g6098), .QN(n5988) );
  SDFFX1 DFF_839_Q_reg ( .D(g29262), .SI(g6098), .SE(test_se), .CLK(CK), .Q(
        g3147), .QN(n5738) );
  SDFFX1 DFF_840_Q_reg ( .D(g24270), .SI(g3147), .SE(test_se), .CLK(CK), .Q(
        g3347), .QN() );
  SDFFX1 DFF_841_Q_reg ( .D(g33581), .SI(g3347), .SE(test_se), .CLK(CK), .Q(
        g2269), .QN(n5410) );
  SDFFX1 DFF_842_Q_reg ( .D(g8358), .SI(g2269), .SE(test_se), .CLK(CK), .Q(
        g191), .QN() );
  SDFFX1 DFF_843_Q_reg ( .D(g24266), .SI(g191), .SE(test_se), .CLK(CK), .Q(
        g2712), .QN() );
  SDFFX1 DFF_844_Q_reg ( .D(g34849), .SI(g2712), .SE(test_se), .CLK(CK), .Q(
        g626), .QN(n5288) );
  SDFFX1 DFF_846_Q_reg ( .D(g33618), .SI(g2729), .SE(test_se), .CLK(CK), .Q(
        g5357), .QN(n5393) );
  SDFFX1 DFF_847_Q_reg ( .D(g34038), .SI(g5357), .SE(test_se), .CLK(CK), .Q(
        test_so58), .QN(n5284) );
  SDFFX1 DFF_848_Q_reg ( .D(g13068), .SI(test_si59), .SE(test_se), .CLK(CK), 
        .Q(g17819), .QN() );
  SDFFX1 DFF_849_Q_reg ( .D(g34032), .SI(g17819), .SE(test_se), .CLK(CK), .Q(
        g4709), .QN(n5518) );
  SDFFX1 DFF_852_Q_reg ( .D(g34803), .SI(g4709), .SE(test_se), .CLK(CK), .Q(
        g2927), .QN() );
  SDFFX1 DFF_853_Q_reg ( .D(g34459), .SI(g2927), .SE(test_se), .CLK(CK), .Q(
        g4340), .QN(n5653) );
  SDFFX1 DFF_854_Q_reg ( .D(g30509), .SI(g4340), .SE(test_se), .CLK(CK), .Q(
        g5929), .QN() );
  SDFFX1 DFF_855_Q_reg ( .D(g34640), .SI(g5929), .SE(test_se), .CLK(CK), .Q(
        g4907), .QN(n5295) );
  SDFFX1 DFF_856_Q_reg ( .D(g14421), .SI(g4907), .SE(test_se), .CLK(CK), .Q(
        g16874), .QN() );
  SDFFX1 DFF_857_Q_reg ( .D(g28069), .SI(g16874), .SE(test_se), .CLK(CK), .Q(
        g4035), .QN() );
  SDFFX1 DFF_858_Q_reg ( .D(g21899), .SI(g4035), .SE(test_se), .CLK(CK), .Q(
        g2946), .QN() );
  SDFFX1 DFF_859_Q_reg ( .D(g31868), .SI(g2946), .SE(test_se), .CLK(CK), .Q(
        g918), .QN(n5673) );
  SDFFX1 DFF_860_Q_reg ( .D(g26938), .SI(g918), .SE(test_se), .CLK(CK), .Q(
        g4082), .QN() );
  SDFFX1 DFF_861_Q_reg ( .D(g25756), .SI(g4082), .SE(test_se), .CLK(CK), .Q(
        g9743), .QN(n5719) );
  SDFFX1 DFF_862_Q_reg ( .D(g30363), .SI(g9743), .SE(test_se), .CLK(CK), .Q(
        test_so59), .QN(n5838) );
  SDFFX1 DFF_863_Q_reg ( .D(g30334), .SI(test_si60), .SE(test_se), .CLK(CK), 
        .Q(g577), .QN(n5294) );
  SDFFX1 DFF_864_Q_reg ( .D(g33970), .SI(g577), .SE(test_se), .CLK(CK), .Q(
        g1620), .QN(n5791) );
  SDFFX1 DFF_865_Q_reg ( .D(g30391), .SI(g1620), .SE(test_se), .CLK(CK), .Q(
        g2831), .QN(g23759) );
  SDFFX1 DFF_866_Q_reg ( .D(g25615), .SI(g2831), .SE(test_se), .CLK(CK), .Q(
        g667), .QN() );
  SDFFX1 DFF_867_Q_reg ( .D(g33540), .SI(g667), .SE(test_se), .CLK(CK), .Q(
        g930), .QN(n5731) );
  SDFFX1 DFF_868_Q_reg ( .D(g30445), .SI(g930), .SE(test_se), .CLK(CK), .Q(
        g3937), .QN() );
  SDFFX1 DFF_870_Q_reg ( .D(g25617), .SI(g3937), .SE(test_se), .CLK(CK), .Q(
        g817), .QN(n5822) );
  SDFFX1 DFF_871_Q_reg ( .D(g24247), .SI(g817), .SE(test_se), .CLK(CK), .Q(
        g1249), .QN() );
  SDFFX1 DFF_872_Q_reg ( .D(g24215), .SI(g1249), .SE(test_se), .CLK(CK), .Q(
        g837), .QN(n5562) );
  SDFFX1 DFF_873_Q_reg ( .D(g14451), .SI(g837), .SE(test_se), .CLK(CK), .Q(
        g16924), .QN() );
  SDFFX1 DFF_874_Q_reg ( .D(g33964), .SI(g16924), .SE(test_se), .CLK(CK), .Q(
        g599), .QN(n5550) );
  SDFFX1 DFF_875_Q_reg ( .D(g25719), .SI(g599), .SE(test_se), .CLK(CK), .Q(
        g5475), .QN(n5425) );
  SDFFX1 DFF_876_Q_reg ( .D(g29228), .SI(g5475), .SE(test_se), .CLK(CK), .Q(
        test_so60), .QN() );
  SDFFX1 DFF_877_Q_reg ( .D(g30514), .SI(test_si61), .SE(test_se), .CLK(CK), 
        .Q(g5949), .QN() );
  SDFFX1 DFF_878_Q_reg ( .D(g33627), .SI(g5949), .SE(test_se), .CLK(CK), .Q(
        g6682), .QN(n5590) );
  SDFFX1 DFF_880_Q_reg ( .D(g24231), .SI(g6682), .SE(test_se), .CLK(CK), .Q(
        g904), .QN() );
  SDFFX1 DFF_881_Q_reg ( .D(g34615), .SI(g904), .SE(test_se), .CLK(CK), .Q(
        g2873), .QN(n5488) );
  SDFFX1 DFF_882_Q_reg ( .D(g30356), .SI(g2873), .SE(test_se), .CLK(CK), .Q(
        g1854), .QN(n5785) );
  SDFFX1 DFF_883_Q_reg ( .D(g25696), .SI(g1854), .SE(test_se), .CLK(CK), .Q(
        g5084), .QN(n5681) );
  SDFFX1 DFF_884_Q_reg ( .D(g30493), .SI(g5084), .SE(test_se), .CLK(CK), .Q(
        g5603), .QN() );
  SDFFX1 DFF_885_Q_reg ( .D(g8917), .SI(g5603), .SE(test_se), .CLK(CK), .Q(
        g8870), .QN(n5726) );
  SDFFX1 DFF_886_Q_reg ( .D(g33594), .SI(g8870), .SE(test_se), .CLK(CK), .Q(
        g2495), .QN(n5522) );
  SDFFX1 DFF_887_Q_reg ( .D(g34009), .SI(g2495), .SE(test_se), .CLK(CK), .Q(
        g2437), .QN(n5789) );
  SDFFX1 DFF_888_Q_reg ( .D(g30365), .SI(g2437), .SE(test_se), .CLK(CK), .Q(
        g2102), .QN(n5666) );
  SDFFX1 DFF_889_Q_reg ( .D(g33004), .SI(g2102), .SE(test_se), .CLK(CK), .Q(
        g2208), .QN() );
  SDFFX1 DFF_890_Q_reg ( .D(g34018), .SI(g2208), .SE(test_se), .CLK(CK), .Q(
        test_so61), .QN(n5684) );
  SDFFX1 DFF_891_Q_reg ( .D(g25685), .SI(test_si62), .SE(test_se), .CLK(CK), 
        .Q(g4064), .QN(n5416) );
  SDFFX1 DFF_892_Q_reg ( .D(g34040), .SI(g4064), .SE(test_se), .CLK(CK), .Q(
        g4899), .QN(n5517) );
  SDFFX1 DFF_893_Q_reg ( .D(g25639), .SI(g4899), .SE(test_se), .CLK(CK), .Q(
        g2719), .QN(n5465) );
  SDFFX1 DFF_894_Q_reg ( .D(g34029), .SI(g2719), .SE(test_se), .CLK(CK), .Q(
        g4785), .QN(n5361) );
  SDFFX1 DFF_895_Q_reg ( .D(g30488), .SI(g4785), .SE(test_se), .CLK(CK), .Q(
        g5583), .QN() );
  SDFFX1 DFF_896_Q_reg ( .D(g34600), .SI(g5583), .SE(test_se), .CLK(CK), .Q(
        g781), .QN(n5551) );
  SDFFX1 DFF_897_Q_reg ( .D(g29300), .SI(g781), .SE(test_se), .CLK(CK), .Q(
        g6173), .QN(n5810) );
  SDFFX1 DFF_898_Q_reg ( .D(g14705), .SI(g6173), .SE(test_se), .CLK(CK), .Q(
        g17743), .QN() );
  SDFFX1 DFF_899_Q_reg ( .D(g34802), .SI(g17743), .SE(test_se), .CLK(CK), .Q(
        g2917), .QN() );
  SDFFX1 DFF_900_Q_reg ( .D(g25614), .SI(g2917), .SE(test_se), .CLK(CK), .Q(
        g686), .QN() );
  SDFFX1 DFF_901_Q_reg ( .D(g28058), .SI(g686), .SE(test_se), .CLK(CK), .Q(
        g1252), .QN(n5554) );
  SDFFX1 DFF_902_Q_reg ( .D(g29225), .SI(g1252), .SE(test_se), .CLK(CK), .Q(
        g671), .QN() );
  SDFFX1 DFF_903_Q_reg ( .D(g33580), .SI(g671), .SE(test_se), .CLK(CK), .Q(
        test_so62), .QN(n5760) );
  SDFFX1 DFF_904_Q_reg ( .D(g30532), .SI(test_si63), .SE(test_se), .CLK(CK), 
        .Q(g6283), .QN() );
  SDFFX1 DFF_905_Q_reg ( .D(g17845), .SI(g6283), .SE(test_se), .CLK(CK), .Q(
        g14705), .QN(n5586) );
  SDFFX1 DFF_906_Q_reg ( .D(g17674), .SI(g14705), .SE(test_se), .CLK(CK), .Q(
        g17519), .QN() );
  SDFFX1 DFF_909_Q_reg ( .D(g8783), .SI(g17519), .SE(test_se), .CLK(CK), .Q(
        g8784), .QN(DFF_909_n1) );
  SDFFX1 DFF_910_Q_reg ( .D(g33054), .SI(g8784), .SE(test_se), .CLK(CK), .Q(
        g5527), .QN(n5389) );
  SDFFX1 DFF_911_Q_reg ( .D(g26962), .SI(g5527), .SE(test_se), .CLK(CK), .Q(
        g4489), .QN() );
  SDFFX1 DFF_912_Q_reg ( .D(g33564), .SI(g4489), .SE(test_se), .CLK(CK), .Q(
        g1974), .QN(n5450) );
  SDFFX1 DFF_913_Q_reg ( .D(g32984), .SI(g1974), .SE(test_se), .CLK(CK), .Q(
        g1270), .QN(n5716) );
  SDFFX1 DFF_914_Q_reg ( .D(g34039), .SI(g1270), .SE(test_se), .CLK(CK), .Q(
        g4966), .QN(n5706) );
  SDFFX1 DFF_916_Q_reg ( .D(g33065), .SI(g4966), .SE(test_se), .CLK(CK), .Q(
        g6227), .QN(n5568) );
  SDFFX1 DFF_917_Q_reg ( .D(g30443), .SI(g6227), .SE(test_se), .CLK(CK), .Q(
        g3929), .QN() );
  SDFFX1 DFF_918_Q_reg ( .D(g29291), .SI(g3929), .SE(test_se), .CLK(CK), .Q(
        g5503), .QN(n5737) );
  SDFFX1 DFF_919_Q_reg ( .D(g24279), .SI(g5503), .SE(test_se), .CLK(CK), .Q(
        test_so63), .QN() );
  SDFFX1 DFF_920_Q_reg ( .D(g30508), .SI(test_si64), .SE(test_se), .CLK(CK), 
        .Q(g5925), .QN() );
  SDFFX1 DFF_921_Q_reg ( .D(g29232), .SI(g5925), .SE(test_se), .CLK(CK), .Q(
        g1124), .QN(n5692) );
  SDFFX1 DFF_922_Q_reg ( .D(g34269), .SI(g1124), .SE(test_se), .CLK(CK), .Q(
        g4955), .QN(n5614) );
  SDFFX1 DFF_923_Q_reg ( .D(g30464), .SI(g4955), .SE(test_se), .CLK(CK), .Q(
        g5224), .QN() );
  SDFFX1 DFF_924_Q_reg ( .D(g33988), .SI(g5224), .SE(test_se), .CLK(CK), .Q(
        g2012), .QN(n5790) );
  SDFFX1 DFF_925_Q_reg ( .D(g30522), .SI(g2012), .SE(test_se), .CLK(CK), .Q(
        g6203), .QN(n5574) );
  SDFFX1 DFF_926_Q_reg ( .D(g25708), .SI(g6203), .SE(test_se), .CLK(CK), .Q(
        g5120), .QN() );
  SDFFX1 DFF_927_Q_reg ( .D(g14662), .SI(g5120), .SE(test_se), .CLK(CK), .Q(
        g17674), .QN() );
  SDFFX1 DFF_928_Q_reg ( .D(g30374), .SI(g17674), .SE(test_se), .CLK(CK), .Q(
        g2389), .QN(n5631) );
  SDFFX1 DFF_929_Q_reg ( .D(g26953), .SI(g2389), .SE(test_se), .CLK(CK), .Q(
        g4438), .QN() );
  SDFFX1 DFF_930_Q_reg ( .D(g34008), .SI(g4438), .SE(test_se), .CLK(CK), .Q(
        g2429), .QN(n5814) );
  SDFFX1 DFF_931_Q_reg ( .D(g34444), .SI(g2429), .SE(test_se), .CLK(CK), .Q(
        g2787), .QN(n5610) );
  SDFFX1 DFF_932_Q_reg ( .D(g34731), .SI(g2787), .SE(test_se), .CLK(CK), .Q(
        test_so64), .QN(n5623) );
  SDFFX1 DFF_933_Q_reg ( .D(g33606), .SI(test_si65), .SE(test_se), .CLK(CK), 
        .Q(g2675), .QN(n5457) );
  SDFFX1 DFF_934_Q_reg ( .D(g24334), .SI(g2675), .SE(test_se), .CLK(CK), .Q(
        g29218), .QN(n5541) );
  SDFFX1 DFF_935_Q_reg ( .D(g34265), .SI(g29218), .SE(test_se), .CLK(CK), .Q(
        g4836), .QN(n5713) );
  SDFFX1 DFF_936_Q_reg ( .D(g30340), .SI(g4836), .SE(test_se), .CLK(CK), .Q(
        g1199), .QN() );
  SDFFX1 DFF_937_Q_reg ( .D(g24257), .SI(g1199), .SE(test_se), .CLK(CK), .Q(
        g19357), .QN(n5401) );
  SDFFX1 DFF_938_Q_reg ( .D(g30482), .SI(g19357), .SE(test_se), .CLK(CK), .Q(
        g5547), .QN() );
  SDFFX1 DFF_941_Q_reg ( .D(g34604), .SI(g5547), .SE(test_se), .CLK(CK), .Q(
        g2138), .QN(n5275) );
  SDFFX1 DFF_942_Q_reg ( .D(g13926), .SI(g2138), .SE(test_se), .CLK(CK), .Q(
        g16744), .QN() );
  SDFFX1 DFF_943_Q_reg ( .D(g33591), .SI(g16744), .SE(test_se), .CLK(CK), .Q(
        g2338), .QN(n5310) );
  SDFFX1 DFF_944_Q_reg ( .D(g8918), .SI(g2338), .SE(test_se), .CLK(CK), .Q(
        g8919), .QN(DFF_944_n1) );
  SDFFX1 DFF_945_Q_reg ( .D(g30525), .SI(g8919), .SE(test_se), .CLK(CK), .Q(
        g6247), .QN() );
  SDFFX1 DFF_946_Q_reg ( .D(g26929), .SI(g6247), .SE(test_se), .CLK(CK), .Q(
        g2791), .QN() );
  SDFFX1 DFF_947_Q_reg ( .D(g30448), .SI(g2791), .SE(test_se), .CLK(CK), .Q(
        test_so65), .QN() );
  SDFFX1 DFF_948_Q_reg ( .D(g34602), .SI(test_si66), .SE(test_se), .CLK(CK), 
        .Q(g1291), .QN(n2549) );
  SDFFX1 DFF_949_Q_reg ( .D(g30513), .SI(g1291), .SE(test_se), .CLK(CK), .Q(
        g5945), .QN() );
  SDFFX1 DFF_950_Q_reg ( .D(g30469), .SI(g5945), .SE(test_se), .CLK(CK), .Q(
        g5244), .QN() );
  SDFFX1 DFF_951_Q_reg ( .D(g33608), .SI(g5244), .SE(test_se), .CLK(CK), .Q(
        g2759), .QN() );
  SDFFX1 DFF_952_Q_reg ( .D(g33626), .SI(g2759), .SE(test_se), .CLK(CK), .Q(
        g6741), .QN(n5398) );
  SDFFX1 DFF_953_Q_reg ( .D(g34725), .SI(g6741), .SE(test_se), .CLK(CK), .Q(
        g785), .QN(n5293) );
  SDFFX1 DFF_954_Q_reg ( .D(g30342), .SI(g785), .SE(test_se), .CLK(CK), .Q(
        g1259), .QN(n5553) );
  SDFFX1 DFF_955_Q_reg ( .D(g29267), .SI(g1259), .SE(test_se), .CLK(CK), .Q(
        g3484), .QN(n5668) );
  SDFFX1 DFF_956_Q_reg ( .D(g25593), .SI(g3484), .SE(test_se), .CLK(CK), .Q(
        g209), .QN(n5595) );
  SDFFX1 DFF_957_Q_reg ( .D(g30548), .SI(g209), .SE(test_se), .CLK(CK), .Q(
        g6609), .QN() );
  SDFFX1 DFF_958_Q_reg ( .D(g33052), .SI(g6609), .SE(test_se), .CLK(CK), .Q(
        g5517), .QN() );
  SDFFX1 DFF_959_Q_reg ( .D(g34012), .SI(g5517), .SE(test_se), .CLK(CK), .Q(
        g2449), .QN(n5798) );
  SDFFX1 DFF_960_Q_reg ( .D(g34017), .SI(g2449), .SE(test_se), .CLK(CK), .Q(
        test_so66), .QN(n5858) );
  SDFFX1 DFF_961_Q_reg ( .D(g29218), .SI(test_si67), .SE(test_se), .CLK(CK), 
        .Q(n9281), .QN(DFF_961_n1) );
  SDFFX1 DFF_962_Q_reg ( .D(g24263), .SI(n9281), .SE(test_se), .CLK(CK), .Q(
        g2715), .QN(n5299) );
  SDFFX1 DFF_963_Q_reg ( .D(g26912), .SI(g2715), .SE(test_se), .CLK(CK), .Q(
        g936), .QN(n5557) );
  SDFFX1 DFF_964_Q_reg ( .D(g30364), .SI(g936), .SE(test_se), .CLK(CK), .Q(
        g2098), .QN(n5280) );
  SDFFX1 DFF_965_Q_reg ( .D(g34254), .SI(g2098), .SE(test_se), .CLK(CK), .Q(
        g4462), .QN(n5671) );
  SDFFX1 DFF_966_Q_reg ( .D(g34251), .SI(g4462), .SE(test_se), .CLK(CK), .Q(
        g604), .QN(n5473) );
  SDFFX1 DFF_967_Q_reg ( .D(g30560), .SI(g604), .SE(test_se), .CLK(CK), .Q(
        g6589), .QN() );
  SDFFX1 DFF_968_Q_reg ( .D(g33983), .SI(g6589), .SE(test_se), .CLK(CK), .Q(
        n9280), .QN(n5686) );
  SDFFX1 DFF_970_Q_reg ( .D(g13085), .SI(n9280), .SE(test_se), .CLK(CK), .Q(
        g17845), .QN() );
  SDFFX1 DFF_971_Q_reg ( .D(g13099), .SI(g17845), .SE(test_se), .CLK(CK), .Q(
        g17871), .QN() );
  SDFFX1 DFF_972_Q_reg ( .D(g24204), .SI(g17871), .SE(test_se), .CLK(CK), .Q(
        g429), .QN() );
  SDFFX1 DFF_973_Q_reg ( .D(g33980), .SI(g429), .SE(test_se), .CLK(CK), .Q(
        g1870), .QN(n5813) );
  SDFFX1 DFF_974_Q_reg ( .D(g34631), .SI(g1870), .SE(test_se), .CLK(CK), .Q(
        test_so67), .QN(n5638) );
  SDFFX1 DFF_977_Q_reg ( .D(g29243), .SI(test_si68), .SE(test_se), .CLK(CK), 
        .Q(g1825), .QN() );
  SDFFX1 DFF_979_Q_reg ( .D(g25623), .SI(g1825), .SE(test_se), .CLK(CK), .Q(
        g1008), .QN(n5321) );
  SDFFX1 DFF_980_Q_reg ( .D(g26950), .SI(g1008), .SE(test_se), .CLK(CK), .Q(
        g4392), .QN(n5710) );
  SDFFX1 DFF_981_Q_reg ( .D(g8178), .SI(g4392), .SE(test_se), .CLK(CK), .Q(
        g8283), .QN() );
  SDFFX1 DFF_982_Q_reg ( .D(g30431), .SI(g8283), .SE(test_se), .CLK(CK), .Q(
        g3546), .QN() );
  SDFFX1 DFF_983_Q_reg ( .D(g30467), .SI(g3546), .SE(test_se), .CLK(CK), .Q(
        g5236), .QN() );
  SDFFX1 DFF_984_Q_reg ( .D(g30353), .SI(g5236), .SE(test_se), .CLK(CK), .Q(
        g1768), .QN(n5834) );
  SDFFX1 DFF_985_Q_reg ( .D(g34467), .SI(g1768), .SE(test_se), .CLK(CK), .Q(
        g4854), .QN() );
  SDFFX1 DFF_986_Q_reg ( .D(g30442), .SI(g4854), .SE(test_se), .CLK(CK), .Q(
        g3925), .QN() );
  SDFFX1 DFF_987_Q_reg ( .D(g29305), .SI(g3925), .SE(test_se), .CLK(CK), .Q(
        g6509), .QN() );
  SDFFX1 DFF_988_Q_reg ( .D(g25616), .SI(g6509), .SE(test_se), .CLK(CK), .Q(
        g732), .QN(n5732) );
  SDFFX1 DFF_989_Q_reg ( .D(g29252), .SI(g732), .SE(test_se), .CLK(CK), .Q(
        g2504), .QN() );
  SDFFX1 DFF_990_Q_reg ( .D(g13272), .SI(g2504), .SE(test_se), .CLK(CK), .Q(
        test_so68), .QN(n5319) );
  SDFFX1 DFF_991_Q_reg ( .D(g4519), .SI(test_si69), .SE(test_se), .CLK(CK), 
        .Q(g4520), .QN() );
  SDFFX1 DFF_992_Q_reg ( .D(g8916), .SI(g4520), .SE(test_se), .CLK(CK), .Q(
        g8917), .QN(DFF_992_n1) );
  SDFFX1 DFF_993_Q_reg ( .D(g33003), .SI(g8917), .SE(test_se), .CLK(CK), .Q(
        g2185), .QN(n5376) );
  SDFFX1 DFF_994_Q_reg ( .D(g34613), .SI(g2185), .SE(test_se), .CLK(CK), .Q(
        g37), .QN(g23002) );
  SDFFX1 DFF_995_Q_reg ( .D(g16748), .SI(g37), .SE(test_se), .CLK(CK), .Q(
        g4031), .QN() );
  SDFFX1 DFF_996_Q_reg ( .D(g33570), .SI(g4031), .SE(test_se), .CLK(CK), .Q(
        g2070), .QN(n5535) );
  SDFFX1 DFF_997_Q_reg ( .D(g8132), .SI(g2070), .SE(test_se), .CLK(CK), .Q(
        g8235), .QN() );
  SDFFX1 DFF_1000_Q_reg ( .D(g34734), .SI(g8235), .SE(test_se), .CLK(CK), .Q(
        g4176), .QN(n5494) );
  SDFFX1 DFF_1001_Q_reg ( .D(g24275), .SI(g4176), .SE(test_se), .CLK(CK), .Q(
        g11418), .QN(n5435) );
  SDFFX1 DFF_1002_Q_reg ( .D(g7243), .SI(g11418), .SE(test_se), .CLK(CK), .Q(
        g4405), .QN() );
  SDFFX1 DFF_1003_Q_reg ( .D(g14167), .SI(g4405), .SE(test_se), .CLK(CK), .Q(
        g872), .QN() );
  SDFFX1 DFF_1004_Q_reg ( .D(g29302), .SI(g872), .SE(test_se), .CLK(CK), .Q(
        g6181), .QN(n5667) );
  SDFFX1 DFF_1005_Q_reg ( .D(g24349), .SI(g6181), .SE(test_se), .CLK(CK), .Q(
        test_so69), .QN(n5533) );
  SDFFX1 DFF_1006_Q_reg ( .D(g34264), .SI(test_si70), .SE(test_se), .CLK(CK), 
        .Q(g4765), .QN(n5613) );
  SDFFX1 DFF_1007_Q_reg ( .D(g30484), .SI(g4765), .SE(test_se), .CLK(CK), .Q(
        g5563), .QN() );
  SDFFX1 DFF_1008_Q_reg ( .D(g25634), .SI(g5563), .SE(test_se), .CLK(CK), .Q(
        g1395), .QN() );
  SDFFX1 DFF_1009_Q_reg ( .D(g33567), .SI(g1395), .SE(test_se), .CLK(CK), .Q(
        g1913), .QN(n5828) );
  SDFFX1 DFF_1010_Q_reg ( .D(g33585), .SI(g1913), .SE(test_se), .CLK(CK), .Q(
        g2331), .QN(n5513) );
  SDFFX1 DFF_1011_Q_reg ( .D(g30527), .SI(g2331), .SE(test_se), .CLK(CK), .Q(
        g6263), .QN() );
  SDFFX1 DFF_1012_Q_reg ( .D(g34978), .SI(g6263), .SE(test_se), .CLK(CK), .Q(
        n9276), .QN(DFF_1012_n1) );
  SDFFX1 DFF_1013_Q_reg ( .D(g30447), .SI(n9276), .SE(test_se), .CLK(CK), .Q(
        g3945), .QN() );
  SDFFX1 DFF_1014_Q_reg ( .D(g7540), .SI(g3945), .SE(test_se), .CLK(CK), .Q(
        g347), .QN(n5860) );
  SDFFX1 DFF_1016_Q_reg ( .D(g34256), .SI(g347), .SE(test_se), .CLK(CK), .Q(
        g4473), .QN() );
  SDFFX1 DFF_1017_Q_reg ( .D(g25630), .SI(g4473), .SE(test_se), .CLK(CK), .Q(
        g1266), .QN() );
  SDFFX1 DFF_1018_Q_reg ( .D(g29290), .SI(g1266), .SE(test_se), .CLK(CK), .Q(
        g5489), .QN(n5660) );
  SDFFX1 DFF_1019_Q_reg ( .D(g29227), .SI(g5489), .SE(test_se), .CLK(CK), .Q(
        test_so70), .QN() );
  SDFFX1 DFF_1020_Q_reg ( .D(g31872), .SI(test_si71), .SE(test_se), .CLK(CK), 
        .Q(g2748), .QN(n5516) );
  SDFFX1 DFF_1021_Q_reg ( .D(g29287), .SI(g2748), .SE(test_se), .CLK(CK), .Q(
        g5471), .QN() );
  SDFFX1 DFF_1022_Q_reg ( .D(g31897), .SI(g5471), .SE(test_se), .CLK(CK), .Q(
        g4540), .QN() );
  SDFFX1 DFF_1023_Q_reg ( .D(g17764), .SI(g4540), .SE(test_se), .CLK(CK), .Q(
        g6723), .QN() );
  SDFFX1 DFF_1024_Q_reg ( .D(g30562), .SI(g6723), .SE(test_se), .CLK(CK), .Q(
        g6605), .QN() );
  SDFFX1 DFF_1025_Q_reg ( .D(g34011), .SI(g6605), .SE(test_se), .CLK(CK), .Q(
        n9274), .QN(n5685) );
  SDFFX1 DFF_1026_Q_reg ( .D(g33996), .SI(n9274), .SE(test_se), .CLK(CK), .Q(
        g2173), .QN(n5857) );
  SDFFX1 DFF_1027_Q_reg ( .D(g21898), .SI(g2173), .SE(test_se), .CLK(CK), .Q(
        g9019), .QN() );
  SDFFX1 DFF_1028_Q_reg ( .D(g33014), .SI(g9019), .SE(test_se), .CLK(CK), .Q(
        g2491), .QN(n5405) );
  SDFFX1 DFF_1029_Q_reg ( .D(g34465), .SI(g2491), .SE(test_se), .CLK(CK), .Q(
        g4849), .QN() );
  SDFFX1 DFF_1030_Q_reg ( .D(g33995), .SI(g4849), .SE(test_se), .CLK(CK), .Q(
        g2169), .QN(n5788) );
  SDFFX1 DFF_1031_Q_reg ( .D(g30372), .SI(g2169), .SE(test_se), .CLK(CK), .Q(
        n9273), .QN(n5624) );
  SDFFX1 DFF_1032_Q_reg ( .D(g30545), .SI(n9273), .SE(test_se), .CLK(CK), .Q(
        test_so71), .QN() );
  SDFFX1 DFF_1033_Q_reg ( .D(g30389), .SI(test_si72), .SE(test_se), .CLK(CK), 
        .Q(g20654), .QN() );
  SDFFX1 DFF_1034_Q_reg ( .D(g33590), .SI(g20654), .SE(test_se), .CLK(CK), .Q(
        g2407), .QN(n5459) );
  SDFFX1 DFF_1035_Q_reg ( .D(g34616), .SI(g2407), .SE(test_se), .CLK(CK), .Q(
        g2868), .QN() );
  SDFFX1 DFF_1036_Q_reg ( .D(g26927), .SI(g2868), .SE(test_se), .CLK(CK), .Q(
        g2767), .QN() );
  SDFFX1 DFF_1037_Q_reg ( .D(g32992), .SI(g2767), .SE(test_se), .CLK(CK), .Q(
        g1783), .QN(n5596) );
  SDFFX1 DFF_1038_Q_reg ( .D(g13895), .SI(g1783), .SE(test_se), .CLK(CK), .Q(
        g16718), .QN() );
  SDFFX1 DFF_1039_Q_reg ( .D(g25631), .SI(g16718), .SE(test_se), .CLK(CK), .Q(
        g1312), .QN(n5466) );
  SDFFX1 DFF_1040_Q_reg ( .D(g30477), .SI(g1312), .SE(test_se), .CLK(CK), .Q(
        g5212), .QN() );
  SDFFX1 DFF_1041_Q_reg ( .D(g34632), .SI(g5212), .SE(test_se), .CLK(CK), .Q(
        g4245), .QN(n5640) );
  SDFFX1 DFF_1042_Q_reg ( .D(g28046), .SI(g4245), .SE(test_se), .CLK(CK), .Q(
        g645), .QN() );
  SDFFX1 DFF_1043_Q_reg ( .D(g9019), .SI(g645), .SE(test_se), .CLK(CK), .Q(
        g4291), .QN() );
  SDFFX1 DFF_1044_Q_reg ( .D(g26896), .SI(g4291), .SE(test_se), .CLK(CK), .Q(
        g20899), .QN(n5657) );
  SDFFX1 DFF_1045_Q_reg ( .D(g25602), .SI(g20899), .SE(test_se), .CLK(CK), .Q(
        test_so72), .QN(n5306) );
  SDFFX1 DFF_1046_Q_reg ( .D(g26916), .SI(test_si73), .SE(test_se), .CLK(CK), 
        .Q(g1129), .QN(n5329) );
  SDFFX1 DFF_1047_Q_reg ( .D(g33578), .SI(g1129), .SE(test_se), .CLK(CK), .Q(
        g2227), .QN(n5538) );
  SDFFX1 DFF_1049_Q_reg ( .D(g8787), .SI(g2227), .SE(test_se), .CLK(CK), .Q(
        g8788), .QN() );
  SDFFX1 DFF_1050_Q_reg ( .D(g33579), .SI(g8788), .SE(test_se), .CLK(CK), .Q(
        g2246), .QN() );
  SDFFX1 DFF_1051_Q_reg ( .D(g30354), .SI(g2246), .SE(test_se), .CLK(CK), .Q(
        g1830), .QN(n5413) );
  SDFFX1 DFF_1052_Q_reg ( .D(g30425), .SI(g1830), .SE(test_se), .CLK(CK), .Q(
        g3590), .QN() );
  SDFFX1 DFF_1053_Q_reg ( .D(g24200), .SI(g3590), .SE(test_se), .CLK(CK), .Q(
        g392), .QN() );
  SDFFX1 DFF_1054_Q_reg ( .D(g33544), .SI(g392), .SE(test_se), .CLK(CK), .Q(
        g1592), .QN(n5362) );
  SDFFX1 DFF_1055_Q_reg ( .D(g25764), .SI(g1592), .SE(test_se), .CLK(CK), .Q(
        g6505), .QN() );
  SDFFX1 DFF_1057_Q_reg ( .D(g24246), .SI(g6505), .SE(test_se), .CLK(CK), .Q(
        g1221), .QN() );
  SDFFX1 DFF_1058_Q_reg ( .D(g30507), .SI(g1221), .SE(test_se), .CLK(CK), .Q(
        g5921), .QN() );
  SDFFX1 DFF_1059_Q_reg ( .D(g26889), .SI(g5921), .SE(test_se), .CLK(CK), .Q(
        g21176), .QN() );
  SDFFX1 DFF_1060_Q_reg ( .D(g30333), .SI(g21176), .SE(test_se), .CLK(CK), .Q(
        test_so73), .QN() );
  SDFFX1 DFF_1061_Q_reg ( .D(g8291), .SI(test_si74), .SE(test_se), .CLK(CK), 
        .Q(g218), .QN() );
  SDFFX1 DFF_1063_Q_reg ( .D(g32998), .SI(g218), .SE(test_se), .CLK(CK), .Q(
        g1932), .QN(n5829) );
  SDFFX1 DFF_1064_Q_reg ( .D(g32987), .SI(g1932), .SE(test_se), .CLK(CK), .Q(
        g1624), .QN(n5370) );
  SDFFX1 DFF_1065_Q_reg ( .D(g25702), .SI(g1624), .SE(test_se), .CLK(CK), .Q(
        g5062), .QN() );
  SDFFX1 DFF_1066_Q_reg ( .D(g29286), .SI(g5062), .SE(test_se), .CLK(CK), .Q(
        g5462), .QN(n5744) );
  SDFFX1 DFF_1067_Q_reg ( .D(g34606), .SI(g5462), .SE(test_se), .CLK(CK), .Q(
        g2689), .QN(n5347) );
  SDFFX1 DFF_1068_Q_reg ( .D(g33070), .SI(g2689), .SE(test_se), .CLK(CK), .Q(
        g6573), .QN(n5563) );
  SDFFX1 DFF_1069_Q_reg ( .D(g29240), .SI(g6573), .SE(test_se), .CLK(CK), .Q(
        g1677), .QN() );
  SDFFX1 DFF_1070_Q_reg ( .D(g32999), .SI(g1677), .SE(test_se), .CLK(CK), .Q(
        g2028), .QN(n5371) );
  SDFFX1 DFF_1071_Q_reg ( .D(g33605), .SI(g2028), .SE(test_se), .CLK(CK), .Q(
        g2671), .QN(n5278) );
  SDFFX1 DFF_1072_Q_reg ( .D(g24255), .SI(g2671), .SE(test_se), .CLK(CK), .Q(
        g10527), .QN() );
  SDFFX1 DFF_1073_Q_reg ( .D(g26945), .SI(g10527), .SE(test_se), .CLK(CK), .Q(
        g7243), .QN() );
  SDFFX1 DFF_1074_Q_reg ( .D(n1278), .SI(g7243), .SE(test_se), .CLK(CK), .Q(
        test_so74), .QN(n5325) );
  SDFFX1 DFF_1075_Q_reg ( .D(g33558), .SI(test_si75), .SE(test_se), .CLK(CK), 
        .Q(g1848), .QN(n5464) );
  SDFFX1 DFF_1078_Q_reg ( .D(g25699), .SI(g1848), .SE(test_se), .CLK(CK), .Q(
        g20557), .QN(n5669) );
  SDFFX1 DFF_1079_Q_reg ( .D(g29289), .SI(g20557), .SE(test_se), .CLK(CK), .Q(
        g5485), .QN(n5869) );
  SDFFX1 DFF_1080_Q_reg ( .D(g30388), .SI(g5485), .SE(test_se), .CLK(CK), .Q(
        g2741), .QN(n5349) );
  SDFFX1 DFF_1081_Q_reg ( .D(g12184), .SI(g2741), .SE(test_se), .CLK(CK), .Q(
        g11678), .QN(n5482) );
  SDFFX1 DFF_1082_Q_reg ( .D(g29254), .SI(g11678), .SE(test_se), .CLK(CK), .Q(
        g2638), .QN() );
  SDFFX1 DFF_1083_Q_reg ( .D(g28074), .SI(g2638), .SE(test_se), .CLK(CK), .Q(
        g4122), .QN() );
  SDFFX1 DFF_1084_Q_reg ( .D(g34450), .SI(g4122), .SE(test_se), .CLK(CK), .Q(
        g4322), .QN(n5506) );
  SDFFX1 DFF_1085_Q_reg ( .D(g30512), .SI(g4322), .SE(test_se), .CLK(CK), .Q(
        g5941), .QN() );
  SDFFX1 DFF_1086_Q_reg ( .D(g33572), .SI(g5941), .SE(test_se), .CLK(CK), .Q(
        g2108), .QN(n5452) );
  SDFFX1 DFF_1087_Q_reg ( .D(g17646), .SI(g2108), .SE(test_se), .CLK(CK), .Q(
        g13068), .QN() );
  SDFFX1 DFF_1088_Q_reg ( .D(g25), .SI(g13068), .SE(test_se), .CLK(CK), .Q(g25), .QN() );
  SDFFX1 DFF_1089_Q_reg ( .D(g33551), .SI(g25), .SE(test_se), .CLK(CK), .Q(
        test_so75), .QN(n5621) );
  SDFFX1 DFF_1090_Q_reg ( .D(g33538), .SI(test_si76), .SE(test_se), .CLK(CK), 
        .Q(g595), .QN(n5476) );
  SDFFX1 DFF_1091_Q_reg ( .D(g33005), .SI(g595), .SE(test_se), .CLK(CK), .Q(
        g2217), .QN(n5512) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24248), .SI(g2217), .SE(test_se), .CLK(CK), .Q(
        n9267), .QN(DFF_1092_n1) );
  SDFFX1 DFF_1093_Q_reg ( .D(g33002), .SI(n9267), .SE(test_se), .CLK(CK), .Q(
        g2066), .QN(n5832) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24234), .SI(g2066), .SE(test_se), .CLK(CK), .Q(
        g1152), .QN(n5618) );
  SDFFX1 DFF_1095_Q_reg ( .D(g30471), .SI(g1152), .SE(test_se), .CLK(CK), .Q(
        g5252), .QN() );
  SDFFX1 DFF_1096_Q_reg ( .D(g34000), .SI(g5252), .SE(test_se), .CLK(CK), .Q(
        g2165), .QN() );
  SDFFX1 DFF_1097_Q_reg ( .D(g34016), .SI(g2165), .SE(test_se), .CLK(CK), .Q(
        g2571), .QN(n5787) );
  SDFFX1 DFF_1098_Q_reg ( .D(g33048), .SI(g2571), .SE(test_se), .CLK(CK), .Q(
        g5176), .QN(n5650) );
  SDFFX1 DFF_1100_Q_reg ( .D(g8283), .SI(g5176), .SE(test_se), .CLK(CK), .Q(
        g8403), .QN() );
  SDFFX1 DFF_1102_Q_reg ( .D(g17819), .SI(g8403), .SE(test_se), .CLK(CK), .Q(
        g14673), .QN(n5581) );
  SDFFX1 DFF_1103_Q_reg ( .D(g25628), .SI(g14673), .SE(test_se), .CLK(CK), .Q(
        test_so76), .QN(n5767) );
  SDFFX1 DFF_1104_Q_reg ( .D(g26934), .SI(test_si77), .SE(test_se), .CLK(CK), 
        .Q(g2827), .QN() );
  SDFFX1 DFF_1106_Q_reg ( .D(g14201), .SI(g2827), .SE(test_se), .CLK(CK), .Q(
        g14217), .QN() );
  SDFFX1 DFF_1107_Q_reg ( .D(g34468), .SI(g14217), .SE(test_se), .CLK(CK), .Q(
        g4859), .QN() );
  SDFFX1 DFF_1108_Q_reg ( .D(g24202), .SI(g4859), .SE(test_se), .CLK(CK), .Q(
        g424), .QN() );
  SDFFX1 DFF_1109_Q_reg ( .D(g33542), .SI(g424), .SE(test_se), .CLK(CK), .Q(
        g1274), .QN(n5730) );
  SDFFX1 DFF_1110_Q_reg ( .D(g17404), .SI(g1274), .SE(test_se), .CLK(CK), .Q(
        g17423), .QN() );
  SDFFX1 DFF_1111_Q_reg ( .D(g33435), .SI(g17423), .SE(test_se), .CLK(CK), .Q(
        n9265), .QN(n6006) );
  SDFFX1 DFF_1112_Q_reg ( .D(g34445), .SI(n9265), .SE(test_se), .CLK(CK), .Q(
        g2803), .QN(n5545) );
  SDFFX1 DFF_1114_Q_reg ( .D(g33555), .SI(g2803), .SE(test_se), .CLK(CK), .Q(
        g1821), .QN() );
  SDFFX1 DFF_1115_Q_reg ( .D(g34013), .SI(g1821), .SE(test_se), .CLK(CK), .Q(
        g2509), .QN() );
  SDFFX1 DFF_1116_Q_reg ( .D(g28091), .SI(g2509), .SE(test_se), .CLK(CK), .Q(
        g5073), .QN() );
  SDFFX1 DFF_1117_Q_reg ( .D(g26919), .SI(g5073), .SE(test_se), .CLK(CK), .Q(
        test_so77), .QN(n5556) );
  SDFFX1 DFF_1118_Q_reg ( .D(g8235), .SI(test_si78), .SE(test_se), .CLK(CK), 
        .Q(g8353), .QN() );
  SDFFX1 DFF_1119_Q_reg ( .D(g17685), .SI(g8353), .SE(test_se), .CLK(CK), .Q(
        g13085), .QN() );
  SDFFX1 DFF_1120_Q_reg ( .D(g30554), .SI(g13085), .SE(test_se), .CLK(CK), .Q(
        g6633), .QN() );
  SDFFX1 DFF_1121_Q_reg ( .D(g29281), .SI(g6633), .SE(test_se), .CLK(CK), .Q(
        g5124), .QN() );
  SDFFX1 DFF_1122_Q_reg ( .D(g17316), .SI(g5124), .SE(test_se), .CLK(CK), .Q(
        g17400), .QN() );
  SDFFX1 DFF_1123_Q_reg ( .D(g30537), .SI(g17400), .SE(test_se), .CLK(CK), .Q(
        g6303), .QN() );
  SDFFX1 DFF_1124_Q_reg ( .D(g28092), .SI(g6303), .SE(test_se), .CLK(CK), .Q(
        g5069), .QN() );
  SDFFX1 DFF_1125_Q_reg ( .D(g34732), .SI(g5069), .SE(test_se), .CLK(CK), .Q(
        g2994), .QN(n5634) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28049), .SI(g2994), .SE(test_se), .CLK(CK), .Q(
        g650), .QN() );
  SDFFX1 DFF_1127_Q_reg ( .D(g33545), .SI(g650), .SE(test_se), .CLK(CK), .Q(
        g1636), .QN(n5549) );
  SDFFX1 DFF_1128_Q_reg ( .D(g30441), .SI(g1636), .SE(test_se), .CLK(CK), .Q(
        g3921), .QN() );
  SDFFX1 DFF_1129_Q_reg ( .D(g29247), .SI(g3921), .SE(test_se), .CLK(CK), .Q(
        test_so78), .QN() );
  SDFFX1 DFF_1130_Q_reg ( .D(g24354), .SI(test_si79), .SE(test_se), .CLK(CK), 
        .Q(g6732), .QN() );
  SDFFX1 DFF_1131_Q_reg ( .D(g25636), .SI(g6732), .SE(test_se), .CLK(CK), .Q(
        g1306), .QN(n5796) );
  SDFFX1 DFF_1133_Q_reg ( .D(g26914), .SI(g1306), .SE(test_se), .CLK(CK), .Q(
        g1061), .QN() );
  SDFFX1 DFF_1134_Q_reg ( .D(g25670), .SI(g1061), .SE(test_se), .CLK(CK), .Q(
        g3462), .QN() );
  SDFFX1 DFF_1135_Q_reg ( .D(g33998), .SI(g3462), .SE(test_se), .CLK(CK), .Q(
        g2181), .QN(n5803) );
  SDFFX1 DFF_1136_Q_reg ( .D(g25626), .SI(g2181), .SE(test_se), .CLK(CK), .Q(
        g956), .QN(n5341) );
  SDFFX1 DFF_1137_Q_reg ( .D(g33977), .SI(g956), .SE(test_se), .CLK(CK), .Q(
        g1756), .QN(n5804) );
  SDFFX1 DFF_1138_Q_reg ( .D(g29297), .SI(g1756), .SE(test_se), .CLK(CK), .Q(
        g5849), .QN(n5736) );
  SDFFX1 DFF_1139_Q_reg ( .D(g28071), .SI(g5849), .SE(test_se), .CLK(CK), .Q(
        g4112), .QN() );
  SDFFX1 DFF_1140_Q_reg ( .D(g30387), .SI(g4112), .SE(test_se), .CLK(CK), .Q(
        n9262), .QN(n5313) );
  SDFFX1 DFF_1141_Q_reg ( .D(g33577), .SI(n9262), .SE(test_se), .CLK(CK), .Q(
        g2197), .QN(n5514) );
  SDFFX1 DFF_1143_Q_reg ( .D(g33592), .SI(g2197), .SE(test_se), .CLK(CK), .Q(
        test_so79), .QN(n5357) );
  SDFFX1 DFF_1144_Q_reg ( .D(g26913), .SI(test_si80), .SE(test_se), .CLK(CK), 
        .Q(g1046), .QN() );
  SDFFX1 DFF_1145_Q_reg ( .D(g28044), .SI(g1046), .SE(test_se), .CLK(CK), .Q(
        g482), .QN(n5820) );
  SDFFX1 DFF_1146_Q_reg ( .D(g26948), .SI(g482), .SE(test_se), .CLK(CK), .Q(
        g4401), .QN() );
  SDFFX1 DFF_1148_Q_reg ( .D(g30344), .SI(g4401), .SE(test_se), .CLK(CK), .Q(
        g1514), .QN(n5364) );
  SDFFX1 DFF_1149_Q_reg ( .D(g26885), .SI(g1514), .SE(test_se), .CLK(CK), .Q(
        g329), .QN(n5766) );
  SDFFX1 DFF_1150_Q_reg ( .D(g33069), .SI(g329), .SE(test_se), .CLK(CK), .Q(
        g6565), .QN(n5386) );
  SDFFX1 DFF_1151_Q_reg ( .D(g34621), .SI(g6565), .SE(test_se), .CLK(CK), .Q(
        g2950), .QN() );
  SDFFX1 DFF_1153_Q_reg ( .D(g28059), .SI(g2950), .SE(test_se), .CLK(CK), .Q(
        g1345), .QN() );
  SDFFX1 DFF_1154_Q_reg ( .D(g25762), .SI(g1345), .SE(test_se), .CLK(CK), .Q(
        g6533), .QN(n5445) );
  SDFFX1 DFF_1155_Q_reg ( .D(g16624), .SI(g6533), .SE(test_se), .CLK(CK), .Q(
        g14421), .QN() );
  SDFFX1 DFF_1157_Q_reg ( .D(g34633), .SI(g14421), .SE(test_se), .CLK(CK), .Q(
        g4727), .QN(n5312) );
  SDFFX1 DFF_1158_Q_reg ( .D(g24352), .SI(g4727), .SE(test_se), .CLK(CK), .Q(
        g12470), .QN(n5434) );
  SDFFX1 DFF_1159_Q_reg ( .D(g26925), .SI(test_si81), .SE(test_se), .CLK(CK), 
        .Q(g1536), .QN() );
  SDFFX1 DFF_1160_Q_reg ( .D(g30446), .SI(g1536), .SE(test_se), .CLK(CK), .Q(
        g3941), .QN() );
  SDFFX1 DFF_1161_Q_reg ( .D(g25597), .SI(g3941), .SE(test_se), .CLK(CK), .Q(
        g370), .QN() );
  SDFFX1 DFF_1162_Q_reg ( .D(g24342), .SI(g370), .SE(test_se), .CLK(CK), .Q(
        g5694), .QN() );
  SDFFX1 DFF_1163_Q_reg ( .D(g30357), .SI(g5694), .SE(test_se), .CLK(CK), .Q(
        g1858), .QN(n5892) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26908), .SI(g1858), .SE(test_se), .CLK(CK), .Q(
        g446), .QN() );
  SDFFX1 DFF_1166_Q_reg ( .D(g30399), .SI(g446), .SE(test_se), .CLK(CK), .Q(
        g3219), .QN() );
  SDFFX1 DFF_1167_Q_reg ( .D(g29242), .SI(g3219), .SE(test_se), .CLK(CK), .Q(
        g1811), .QN() );
  SDFFX1 DFF_1169_Q_reg ( .D(g30547), .SI(g1811), .SE(test_se), .CLK(CK), .Q(
        g6601), .QN() );
  SDFFX1 DFF_1171_Q_reg ( .D(g34010), .SI(g6601), .SE(test_se), .CLK(CK), .Q(
        g2441), .QN(n5856) );
  SDFFX1 DFF_1172_Q_reg ( .D(g33986), .SI(g2441), .SE(test_se), .CLK(CK), .Q(
        g1874), .QN() );
  SDFFX1 DFF_1173_Q_reg ( .D(g34257), .SI(g1874), .SE(test_se), .CLK(CK), .Q(
        test_so81), .QN(n5298) );
  SDFFX1 DFF_1174_Q_reg ( .D(g30544), .SI(test_si82), .SE(test_se), .CLK(CK), 
        .Q(g6581), .QN() );
  SDFFX1 DFF_1175_Q_reg ( .D(g30561), .SI(g6581), .SE(test_se), .CLK(CK), .Q(
        g6597), .QN() );
  SDFFX1 DFF_1176_Q_reg ( .D(g8403), .SI(g6597), .SE(test_se), .CLK(CK), .Q(
        g5008), .QN(n5637) );
  SDFFX1 DFF_1177_Q_reg ( .D(g30430), .SI(g5008), .SE(test_se), .CLK(CK), .Q(
        g3610), .QN() );
  SDFFX1 DFF_1178_Q_reg ( .D(g34799), .SI(g3610), .SE(test_se), .CLK(CK), .Q(
        g2890), .QN() );
  SDFFX1 DFF_1179_Q_reg ( .D(g33565), .SI(g2890), .SE(test_se), .CLK(CK), .Q(
        g1978), .QN(n5845) );
  SDFFX1 DFF_1180_Q_reg ( .D(g33968), .SI(g1978), .SE(test_se), .CLK(CK), .Q(
        g1612), .QN(n5855) );
  SDFFX1 DFF_1181_Q_reg ( .D(g34843), .SI(g1612), .SE(test_se), .CLK(CK), .Q(
        g112), .QN() );
  SDFFX1 DFF_1182_Q_reg ( .D(g34793), .SI(g112), .SE(test_se), .CLK(CK), .Q(
        g2856), .QN() );
  SDFFX1 DFF_1184_Q_reg ( .D(g33566), .SI(g2856), .SE(test_se), .CLK(CK), .Q(
        g1982), .QN(n5462) );
  SDFFX1 DFF_1185_Q_reg ( .D(g17688), .SI(g1982), .SE(test_se), .CLK(CK), .Q(
        g17722), .QN() );
  SDFFX1 DFF_1186_Q_reg ( .D(g30465), .SI(g17722), .SE(test_se), .CLK(CK), .Q(
        test_so82), .QN() );
  SDFFX1 DFF_1187_Q_reg ( .D(g28073), .SI(test_si83), .SE(test_se), .CLK(CK), 
        .Q(g4119), .QN() );
  SDFFX1 DFF_1188_Q_reg ( .D(g24351), .SI(g4119), .SE(test_se), .CLK(CK), .Q(
        g6390), .QN() );
  SDFFX1 DFF_1189_Q_reg ( .D(g30346), .SI(g6390), .SE(test_se), .CLK(CK), .Q(
        g1542), .QN() );
  SDFFX1 DFF_1190_Q_reg ( .D(g21893), .SI(g1542), .SE(test_se), .CLK(CK), .Q(
        g4258), .QN() );
  SDFFX1 DFF_1191_Q_reg ( .D(g8353), .SI(g4258), .SE(test_se), .CLK(CK), .Q(
        g4818), .QN(n5636) );
  SDFFX1 DFF_1192_Q_reg ( .D(g31904), .SI(g4818), .SE(test_se), .CLK(CK), .Q(
        g5033), .QN() );
  SDFFX1 DFF_1193_Q_reg ( .D(g34635), .SI(g5033), .SE(test_se), .CLK(CK), .Q(
        g4717), .QN(n5344) );
  SDFFX1 DFF_1194_Q_reg ( .D(g25637), .SI(g4717), .SE(test_se), .CLK(CK), .Q(
        g1554), .QN(n5768) );
  SDFFX1 DFF_1195_Q_reg ( .D(g29274), .SI(g1554), .SE(test_se), .CLK(CK), .Q(
        g3849), .QN(n5735) );
  SDFFX1 DFF_1196_Q_reg ( .D(g14828), .SI(g3849), .SE(test_se), .CLK(CK), .Q(
        g17778), .QN() );
  SDFFX1 DFF_1197_Q_reg ( .D(g30396), .SI(g17778), .SE(test_se), .CLK(CK), .Q(
        g3199), .QN() );
  SDFFX1 DFF_1198_Q_reg ( .D(g25735), .SI(g3199), .SE(test_se), .CLK(CK), .Q(
        test_so83), .QN(n5887) );
  SDFFX1 DFF_1199_Q_reg ( .D(g34037), .SI(test_si84), .SE(test_se), .CLK(CK), 
        .Q(g4975), .QN(n5360) );
  SDFFX1 DFF_1200_Q_reg ( .D(g34791), .SI(g4975), .SE(test_se), .CLK(CK), .Q(
        g790), .QN(n5292) );
  SDFFX1 DFF_1201_Q_reg ( .D(g30520), .SI(g790), .SE(test_se), .CLK(CK), .Q(
        g5913), .QN() );
  SDFFX1 DFF_1202_Q_reg ( .D(g30358), .SI(g5913), .SE(test_se), .CLK(CK), .Q(
        g1902), .QN(n5837) );
  SDFFX1 DFF_1203_Q_reg ( .D(g29299), .SI(g1902), .SE(test_se), .CLK(CK), .Q(
        g6163), .QN() );
  SDFFX1 DFF_1204_Q_reg ( .D(g25690), .SI(g6163), .SE(test_se), .CLK(CK), .Q(
        g4125), .QN() );
  SDFFX1 DFF_1205_Q_reg ( .D(g28096), .SI(g4125), .SE(test_se), .CLK(CK), .Q(
        g4821), .QN(n5880) );
  SDFFX1 DFF_1206_Q_reg ( .D(g28088), .SI(g4821), .SE(test_se), .CLK(CK), .Q(
        g4939), .QN(n5776) );
  SDFFX1 DFF_1207_Q_reg ( .D(g24241), .SI(g4939), .SE(test_se), .CLK(CK), .Q(
        g19334), .QN(n5392) );
  SDFFX1 DFF_1208_Q_reg ( .D(g30397), .SI(g19334), .SE(test_se), .CLK(CK), .Q(
        g3207), .QN() );
  SDFFX1 DFF_1209_Q_reg ( .D(g4520), .SI(g3207), .SE(test_se), .CLK(CK), .Q(
        g4483), .QN() );
  SDFFX1 DFF_1210_Q_reg ( .D(g30409), .SI(g4483), .SE(test_se), .CLK(CK), .Q(
        test_so84), .QN() );
  SDFFX1 DFF_1211_Q_reg ( .D(g29284), .SI(test_si85), .SE(test_se), .CLK(CK), 
        .Q(g5142), .QN(n5658) );
  SDFFX1 DFF_1212_Q_reg ( .D(g30470), .SI(g5142), .SE(test_se), .CLK(CK), .Q(
        g5248), .QN() );
  SDFFX1 DFF_1213_Q_reg ( .D(g30367), .SI(g5248), .SE(test_se), .CLK(CK), .Q(
        g2126), .QN(n5891) );
  SDFFX1 DFF_1214_Q_reg ( .D(g24273), .SI(g2126), .SE(test_se), .CLK(CK), .Q(
        g3694), .QN() );
  SDFFX1 DFF_1215_Q_reg ( .D(g29288), .SI(g3694), .SE(test_se), .CLK(CK), .Q(
        g5481), .QN(n5805) );
  SDFFX1 DFF_1216_Q_reg ( .D(g30359), .SI(g5481), .SE(test_se), .CLK(CK), .Q(
        g1964), .QN(n5315) );
  SDFFX1 DFF_1217_Q_reg ( .D(g25698), .SI(g1964), .SE(test_se), .CLK(CK), .Q(
        g5097), .QN(n5753) );
  SDFFX1 DFF_1218_Q_reg ( .D(g30398), .SI(g5097), .SE(test_se), .CLK(CK), .Q(
        g3215), .QN() );
  SDFFX1 DFF_1219_Q_reg ( .D(g13906), .SI(g3215), .SE(test_se), .CLK(CK), .Q(
        g16748), .QN() );
  SDFFX1 DFF_1220_Q_reg ( .D(g33079), .SI(g16748), .SE(test_se), .CLK(CK), .Q(
        n9255), .QN(n6005) );
  SDFFX1 DFF_1221_Q_reg ( .D(g26952), .SI(n9255), .SE(test_se), .CLK(CK), .Q(
        g4427), .QN() );
  SDFFX1 DFF_1222_Q_reg ( .D(g34974), .SI(g4427), .SE(test_se), .CLK(CK), .Q(
        test_so85), .QN() );
  SDFFX1 DFF_1223_Q_reg ( .D(g26928), .SI(test_si86), .SE(test_se), .CLK(CK), 
        .Q(g2779), .QN() );
  SDFFX1 DFF_1224_Q_reg ( .D(g8785), .SI(g2779), .SE(test_se), .CLK(CK), .Q(
        g8786), .QN(n5694) );
  SDFFX1 DFF_1225_Q_reg ( .D(g26954), .SI(g8786), .SE(test_se), .CLK(CK), .Q(
        g7245), .QN(DFF_1225_n1) );
  SDFFX1 DFF_1226_Q_reg ( .D(g30351), .SI(g7245), .SE(test_se), .CLK(CK), .Q(
        g1720), .QN(n5780) );
  SDFFX1 DFF_1227_Q_reg ( .D(g31871), .SI(g1720), .SE(test_se), .CLK(CK), .Q(
        g1367), .QN() );
  SDFFX1 DFF_1228_Q_reg ( .D(g9553), .SI(g1367), .SE(test_se), .CLK(CK), .Q(
        g5112), .QN() );
  SDFFX1 DFF_1229_Q_reg ( .D(g34978), .SI(g5112), .SE(test_se), .CLK(CK), .Q(
        g19), .QN() );
  SDFFX1 DFF_1230_Q_reg ( .D(g26939), .SI(g19), .SE(test_se), .CLK(CK), .Q(
        g4145), .QN() );
  SDFFX1 DFF_1231_Q_reg ( .D(g33994), .SI(g4145), .SE(test_se), .CLK(CK), .Q(
        g2161), .QN(n5812) );
  SDFFX1 DFF_1232_Q_reg ( .D(g25596), .SI(g2161), .SE(test_se), .CLK(CK), .Q(
        g376), .QN(n5633) );
  SDFFX1 DFF_1233_Q_reg ( .D(g33586), .SI(g376), .SE(test_se), .CLK(CK), .Q(
        g2361), .QN(n5537) );
  SDFFX1 DFF_1234_Q_reg ( .D(g21901), .SI(g2361), .SE(test_se), .CLK(CK), .Q(
        g11447), .QN(DFF_1234_n1) );
  SDFFX1 DFF_1235_Q_reg ( .D(g31866), .SI(test_si87), .SE(test_se), .CLK(CK), 
        .Q(g582), .QN(n5552) );
  SDFFX1 DFF_1236_Q_reg ( .D(g33000), .SI(g582), .SE(test_se), .CLK(CK), .Q(
        g2051), .QN() );
  SDFFX1 DFF_1237_Q_reg ( .D(g26918), .SI(g2051), .SE(test_se), .CLK(CK), .Q(
        g1193), .QN() );
  SDFFX1 DFF_1240_Q_reg ( .D(g30373), .SI(g1193), .SE(test_se), .CLK(CK), .Q(
        g2327), .QN(n5841) );
  SDFFX1 DFF_1241_Q_reg ( .D(g28056), .SI(g2327), .SE(test_se), .CLK(CK), .Q(
        g907), .QN(n5555) );
  SDFFX1 DFF_1242_Q_reg ( .D(g34601), .SI(g907), .SE(test_se), .CLK(CK), .Q(
        g947), .QN(n5286) );
  SDFFX1 DFF_1243_Q_reg ( .D(g30355), .SI(g947), .SE(test_se), .CLK(CK), .Q(
        g1834), .QN(n5665) );
  SDFFX1 DFF_1244_Q_reg ( .D(g30426), .SI(g1834), .SE(test_se), .CLK(CK), .Q(
        g3594), .QN() );
  SDFFX1 DFF_1245_Q_reg ( .D(g34805), .SI(g3594), .SE(test_se), .CLK(CK), .Q(
        g2999), .QN() );
  SDFFX1 DFF_1247_Q_reg ( .D(g34002), .SI(g2999), .SE(test_se), .CLK(CK), .Q(
        g2303), .QN(n5794) );
  SDFFX1 DFF_1248_Q_reg ( .D(g17778), .SI(g2303), .SE(test_se), .CLK(CK), .Q(
        g17688), .QN() );
  SDFFX1 DFF_1250_Q_reg ( .D(g28053), .SI(g17688), .SE(test_se), .CLK(CK), .Q(
        test_so87), .QN() );
  SDFFX1 DFF_1251_Q_reg ( .D(g29229), .SI(test_si88), .SE(test_se), .CLK(CK), 
        .Q(g723), .QN(n5826) );
  SDFFX1 DFF_1252_Q_reg ( .D(g33620), .SI(g723), .SE(test_se), .CLK(CK), .Q(
        g5703), .QN(n5397) );
  SDFFX1 DFF_1253_Q_reg ( .D(g34722), .SI(g5703), .SE(test_se), .CLK(CK), .Q(
        g546), .QN(n5492) );
  SDFFX1 DFF_1254_Q_reg ( .D(g33599), .SI(g546), .SE(test_se), .CLK(CK), .Q(
        g2472), .QN(n5619) );
  SDFFX1 DFF_1255_Q_reg ( .D(g30515), .SI(g2472), .SE(test_se), .CLK(CK), .Q(
        g5953), .QN() );
  SDFFX1 DFF_1256_Q_reg ( .D(g25649), .SI(g5953), .SE(test_se), .CLK(CK), .Q(
        g8277), .QN() );
  SDFFX1 DFF_1258_Q_reg ( .D(g33979), .SI(g8277), .SE(test_se), .CLK(CK), .Q(
        g1740), .QN() );
  SDFFX1 DFF_1259_Q_reg ( .D(g30417), .SI(g1740), .SE(test_se), .CLK(CK), .Q(
        g3550), .QN() );
  SDFFX1 DFF_1260_Q_reg ( .D(g25683), .SI(g3550), .SE(test_se), .CLK(CK), .Q(
        g3845), .QN(n5886) );
  SDFFX1 DFF_1261_Q_reg ( .D(g33574), .SI(g3845), .SE(test_se), .CLK(CK), .Q(
        g2116), .QN(n5463) );
  SDFFX1 DFF_1262_Q_reg ( .D(g17813), .SI(g2116), .SE(test_se), .CLK(CK), .Q(
        g14635), .QN(n5582) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30410), .SI(g14635), .SE(test_se), .CLK(CK), .Q(
        test_so88), .QN() );
  SDFFX1 DFF_1264_Q_reg ( .D(g30454), .SI(test_si89), .SE(test_se), .CLK(CK), 
        .Q(g3913), .QN() );
  SDFFX1 DFF_1265_Q_reg ( .D(g34024), .SI(g3913), .SE(test_se), .CLK(CK), .Q(
        g10306), .QN() );
  SDFFX1 DFF_1266_Q_reg ( .D(g33547), .SI(g10306), .SE(test_se), .CLK(CK), .Q(
        g1687), .QN() );
  SDFFX1 DFF_1267_Q_reg ( .D(g30386), .SI(g1687), .SE(test_se), .CLK(CK), .Q(
        g2681), .QN(n5777) );
  SDFFX1 DFF_1268_Q_reg ( .D(g33596), .SI(g2681), .SE(test_se), .CLK(CK), .Q(
        g2533), .QN(n5761) );
  SDFFX1 DFF_1269_Q_reg ( .D(g26887), .SI(g2533), .SE(test_se), .CLK(CK), .Q(
        g324), .QN(n5827) );
  SDFFX1 DFF_1270_Q_reg ( .D(g34607), .SI(g324), .SE(test_se), .CLK(CK), .Q(
        g2697), .QN(n5308) );
  SDFFX1 DFF_1272_Q_reg ( .D(g31895), .SI(g2697), .SE(test_se), .CLK(CK), .Q(
        g4417), .QN() );
  SDFFX1 DFF_1273_Q_reg ( .D(g33068), .SI(g4417), .SE(test_se), .CLK(CK), .Q(
        g6561), .QN(n5646) );
  SDFFX1 DFF_1274_Q_reg ( .D(g29233), .SI(g6561), .SE(test_se), .CLK(CK), .Q(
        g1141), .QN(n5691) );
  SDFFX1 DFF_1275_Q_reg ( .D(g24258), .SI(g1141), .SE(test_se), .CLK(CK), .Q(
        g12923), .QN(n5655) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30376), .SI(g12923), .SE(test_se), .CLK(CK), .Q(
        test_so89), .QN(n5779) );
  SDFFX1 DFF_1277_Q_reg ( .D(g33549), .SI(test_si90), .SE(test_se), .CLK(CK), 
        .Q(g1710), .QN(n5412) );
  SDFFX1 DFF_1278_Q_reg ( .D(g29308), .SI(g1710), .SE(test_se), .CLK(CK), .Q(
        g6527), .QN(n5659) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30408), .SI(g6527), .SE(test_se), .CLK(CK), .Q(
        g3255), .QN() );
  SDFFX1 DFF_1281_Q_reg ( .D(g29241), .SI(g3255), .SE(test_se), .CLK(CK), .Q(
        g1691), .QN() );
  SDFFX1 DFF_1282_Q_reg ( .D(g34620), .SI(g1691), .SE(test_se), .CLK(CK), .Q(
        g2936), .QN() );
  SDFFX1 DFF_1283_Q_reg ( .D(g33621), .SI(g2936), .SE(test_se), .CLK(CK), .Q(
        g5644), .QN(n5593) );
  SDFFX1 DFF_1284_Q_reg ( .D(g25707), .SI(g5644), .SE(test_se), .CLK(CK), .Q(
        g5152), .QN(n5883) );
  SDFFX1 DFF_1285_Q_reg ( .D(g24339), .SI(g5152), .SE(test_se), .CLK(CK), .Q(
        g5352), .QN() );
  SDFFX1 DFF_1286_Q_reg ( .D(g11770), .SI(g5352), .SE(test_se), .CLK(CK), .Q(
        g8915), .QN() );
  SDFFX1 DFF_1288_Q_reg ( .D(g34443), .SI(g8915), .SE(test_se), .CLK(CK), .Q(
        g2775), .QN(n5378) );
  SDFFX1 DFF_1289_Q_reg ( .D(g34619), .SI(g2775), .SE(test_se), .CLK(CK), .Q(
        g2922), .QN() );
  SDFFX1 DFF_1290_Q_reg ( .D(g29234), .SI(g2922), .SE(test_se), .CLK(CK), .Q(
        test_so90), .QN(n5864) );
  SDFFX1 DFF_1291_Q_reg ( .D(g30503), .SI(test_si91), .SE(test_se), .CLK(CK), 
        .Q(g5893), .QN() );
  SDFFX1 DFF_1293_Q_reg ( .D(g16718), .SI(g5893), .SE(test_se), .CLK(CK), .Q(
        g16603), .QN() );
  SDFFX1 DFF_1294_Q_reg ( .D(g30550), .SI(g16603), .SE(test_se), .CLK(CK), .Q(
        g6617), .QN() );
  SDFFX1 DFF_1295_Q_reg ( .D(g33001), .SI(g6617), .SE(test_se), .CLK(CK), .Q(
        g2060), .QN(n5507) );
  SDFFX1 DFF_1296_Q_reg ( .D(g33040), .SI(g2060), .SE(test_se), .CLK(CK), .Q(
        g4512), .QN() );
  SDFFX1 DFF_1297_Q_reg ( .D(g30492), .SI(g4512), .SE(test_se), .CLK(CK), .Q(
        g5599), .QN() );
  SDFFX1 DFF_1298_Q_reg ( .D(g25664), .SI(g5599), .SE(test_se), .CLK(CK), .Q(
        g3401), .QN(n5986) );
  SDFFX1 DFF_1299_Q_reg ( .D(g26944), .SI(g3401), .SE(test_se), .CLK(CK), .Q(
        g4366), .QN() );
  SDFFX1 DFF_1300_Q_reg ( .D(g13881), .SI(g4366), .SE(test_se), .CLK(CK), .Q(
        g16722), .QN() );
  SDFFX1 DFF_1301_Q_reg ( .D(g34614), .SI(g16722), .SE(test_se), .CLK(CK), .Q(
        g20652), .QN(n5342) );
  SDFFX1 DFF_1302_Q_reg ( .D(g29260), .SI(g20652), .SE(test_se), .CLK(CK), .Q(
        g3129), .QN(n5861) );
  SDFFX1 DFF_1303_Q_reg ( .D(g16686), .SI(g3129), .SE(test_se), .CLK(CK), .Q(
        test_so91), .QN() );
  SDFFX1 DFF_1304_Q_reg ( .D(g33047), .SI(test_si92), .SE(test_se), .CLK(CK), 
        .Q(g5170), .QN() );
  SDFFX1 DFF_1305_Q_reg ( .D(g24298), .SI(g5170), .SE(test_se), .CLK(CK), .Q(
        g26959), .QN() );
  SDFFX1 DFF_1306_Q_reg ( .D(g25733), .SI(g26959), .SE(test_se), .CLK(CK), .Q(
        g5821), .QN(n5429) );
  SDFFX1 DFF_1307_Q_reg ( .D(g30536), .SI(g5821), .SE(test_se), .CLK(CK), .Q(
        g6299), .QN() );
  SDFFX1 DFF_1308_Q_reg ( .D(n6021), .SI(g6299), .SE(test_se), .CLK(CK), .Q(
        g8416), .QN() );
  SDFFX1 DFF_1310_Q_reg ( .D(g29246), .SI(g8416), .SE(test_se), .CLK(CK), .Q(
        g2079), .QN() );
  SDFFX1 DFF_1311_Q_reg ( .D(g34261), .SI(g2079), .SE(test_se), .CLK(CK), .Q(
        g4698), .QN(n5862) );
  SDFFX1 DFF_1312_Q_reg ( .D(g33611), .SI(g4698), .SE(test_se), .CLK(CK), .Q(
        g3703), .QN(n5399) );
  SDFFX1 DFF_1313_Q_reg ( .D(g25638), .SI(g3703), .SE(test_se), .CLK(CK), .Q(
        g1559), .QN(n5441) );
  SDFFX1 DFF_1314_Q_reg ( .D(g34728), .SI(g1559), .SE(test_se), .CLK(CK), .Q(
        n9247), .QN(n5409) );
  SDFFX1 DFF_1315_Q_reg ( .D(g29222), .SI(n9247), .SE(test_se), .CLK(CK), .Q(
        g411), .QN(n5629) );
  SDFFX1 DFF_1316_Q_reg ( .D(g25742), .SI(g411), .SE(test_se), .CLK(CK), .Q(
        g9682), .QN(n5718) );
  SDFFX1 DFF_1317_Q_reg ( .D(g30449), .SI(test_si93), .SE(test_se), .CLK(CK), 
        .Q(g3953), .QN() );
  SDFFX1 DFF_1319_Q_reg ( .D(g34608), .SI(g3953), .SE(test_se), .CLK(CK), .Q(
        g2704), .QN(n5377) );
  SDFFX1 DFF_1320_Q_reg ( .D(g24345), .SI(g2704), .SE(test_se), .CLK(CK), .Q(
        g6035), .QN(n5528) );
  SDFFX1 DFF_1322_Q_reg ( .D(g34977), .SI(g6035), .SE(test_se), .CLK(CK), .Q(
        n9245), .QN(DFF_1322_n1) );
  SDFFX1 DFF_1323_Q_reg ( .D(g25635), .SI(n9245), .SE(test_se), .CLK(CK), .Q(
        g1300), .QN(n5483) );
  SDFFX1 DFF_1324_Q_reg ( .D(g25686), .SI(g1300), .SE(test_se), .CLK(CK), .Q(
        g4057), .QN(n5711) );
  SDFFX1 DFF_1325_Q_reg ( .D(g30461), .SI(g4057), .SE(test_se), .CLK(CK), .Q(
        g5200), .QN() );
  SDFFX1 DFF_1326_Q_reg ( .D(g34466), .SI(g5200), .SE(test_se), .CLK(CK), .Q(
        g4843), .QN() );
  SDFFX1 DFF_1327_Q_reg ( .D(g31901), .SI(g4843), .SE(test_se), .CLK(CK), .Q(
        g5046), .QN(n5578) );
  SDFFX1 DFF_1328_Q_reg ( .D(g29249), .SI(g5046), .SE(test_se), .CLK(CK), .Q(
        g2250), .QN() );
  SDFFX1 DFF_1329_Q_reg ( .D(g26882), .SI(g2250), .SE(test_se), .CLK(CK), .Q(
        g26885), .QN(n5456) );
  SDFFX1 DFF_1330_Q_reg ( .D(g33041), .SI(g26885), .SE(test_se), .CLK(CK), .Q(
        test_so93), .QN() );
  SDFFX1 DFF_1331_Q_reg ( .D(g33011), .SI(test_si94), .SE(test_se), .CLK(CK), 
        .Q(g2453), .QN(n5373) );
  SDFFX1 DFF_1332_Q_reg ( .D(g25734), .SI(g2453), .SE(test_se), .CLK(CK), .Q(
        g5841), .QN(n5449) );
  SDFFX1 DFF_1335_Q_reg ( .D(g12300), .SI(g5841), .SE(test_se), .CLK(CK), .Q(
        g14694), .QN(n5705) );
  SDFFX1 DFF_1336_Q_reg ( .D(g34618), .SI(g14694), .SE(test_se), .CLK(CK), .Q(
        g2912), .QN() );
  SDFFX1 DFF_1337_Q_reg ( .D(g33010), .SI(g2912), .SE(test_se), .CLK(CK), .Q(
        g2357), .QN(n5276) );
  SDFFX1 DFF_1338_Q_reg ( .D(g8919), .SI(g2357), .SE(test_se), .CLK(CK), .Q(
        g8920), .QN(DFF_1338_n1) );
  SDFFX1 DFF_1339_Q_reg ( .D(g31864), .SI(g8920), .SE(test_se), .CLK(CK), .Q(
        g164), .QN(n5561) );
  SDFFX1 DFF_1340_Q_reg ( .D(g34630), .SI(g164), .SE(test_se), .CLK(CK), .Q(
        g4253), .QN(n5484) );
  SDFFX1 DFF_1341_Q_reg ( .D(g31898), .SI(g4253), .SE(test_se), .CLK(CK), .Q(
        g5016), .QN(n5369) );
  SDFFX1 DFF_1342_Q_reg ( .D(g25653), .SI(g5016), .SE(test_se), .CLK(CK), .Q(
        g3119), .QN(n5423) );
  SDFFX1 DFF_1343_Q_reg ( .D(g25632), .SI(g3119), .SE(test_se), .CLK(CK), .Q(
        g1351), .QN(n5322) );
  SDFFX1 DFF_1344_Q_reg ( .D(g32988), .SI(g1351), .SE(test_se), .CLK(CK), .Q(
        test_so94), .QN() );
  SDFFX1 DFF_1345_Q_reg ( .D(g33616), .SI(test_si95), .SE(test_se), .CLK(CK), 
        .Q(g4519), .QN() );
  SDFFX1 DFF_1346_Q_reg ( .D(g29280), .SI(g4519), .SE(test_se), .CLK(CK), .Q(
        g5115), .QN(n5743) );
  SDFFX1 DFF_1347_Q_reg ( .D(g33609), .SI(g5115), .SE(test_se), .CLK(CK), .Q(
        g3352), .QN(n5604) );
  SDFFX1 DFF_1348_Q_reg ( .D(g30563), .SI(g3352), .SE(test_se), .CLK(CK), .Q(
        g6657), .QN() );
  SDFFX1 DFF_1349_Q_reg ( .D(g33044), .SI(g6657), .SE(test_se), .CLK(CK), .Q(
        g4552), .QN() );
  SDFFX1 DFF_1350_Q_reg ( .D(g30437), .SI(g4552), .SE(test_se), .CLK(CK), .Q(
        g3893), .QN() );
  SDFFX1 DFF_1351_Q_reg ( .D(g30412), .SI(g3893), .SE(test_se), .CLK(CK), .Q(
        g3211), .QN() );
  SDFFX1 DFF_1352_Q_reg ( .D(g17604), .SI(g3211), .SE(test_se), .CLK(CK), .Q(
        g13049), .QN() );
  SDFFX1 DFF_1354_Q_reg ( .D(g16603), .SI(g13049), .SE(test_se), .CLK(CK), .Q(
        g16624), .QN() );
  SDFFX1 DFF_1355_Q_reg ( .D(g30491), .SI(g16624), .SE(test_se), .CLK(CK), .Q(
        g5595), .QN() );
  SDFFX1 DFF_1356_Q_reg ( .D(g30434), .SI(g5595), .SE(test_se), .CLK(CK), .Q(
        g3614), .QN() );
  SDFFX1 DFF_1357_Q_reg ( .D(g34612), .SI(g3614), .SE(test_se), .CLK(CK), .Q(
        test_so95), .QN() );
  SDFFX1 DFF_1358_Q_reg ( .D(g29259), .SI(test_si96), .SE(test_se), .CLK(CK), 
        .Q(g3125), .QN(n5781) );
  SDFFX1 DFF_1359_Q_reg ( .D(g13865), .SI(g3125), .SE(test_se), .CLK(CK), .Q(
        g16686), .QN() );
  SDFFX1 DFF_1360_Q_reg ( .D(g25681), .SI(g16686), .SE(test_se), .CLK(CK), .Q(
        g3821), .QN(n5428) );
  SDFFX1 DFF_1361_Q_reg ( .D(g25687), .SI(g3821), .SE(test_se), .CLK(CK), .Q(
        g4141), .QN(n5612) );
  SDFFX1 DFF_1362_Q_reg ( .D(g33617), .SI(g4141), .SE(test_se), .CLK(CK), .Q(
        g4570), .QN() );
  SDFFX1 DFF_1363_Q_reg ( .D(g30479), .SI(g4570), .SE(test_se), .CLK(CK), .Q(
        g5272), .QN() );
  SDFFX1 DFF_1364_Q_reg ( .D(g29256), .SI(g5272), .SE(test_se), .CLK(CK), .Q(
        g2735), .QN(n5600) );
  SDFFX1 DFF_1365_Q_reg ( .D(g28054), .SI(g2735), .SE(test_se), .CLK(CK), .Q(
        g728), .QN() );
  SDFFX1 DFF_1366_Q_reg ( .D(g30535), .SI(g728), .SE(test_se), .CLK(CK), .Q(
        g6295), .QN() );
  SDFFX1 DFF_1368_Q_reg ( .D(g30385), .SI(g6295), .SE(test_se), .CLK(CK), .Q(
        g2661), .QN(n5418) );
  SDFFX1 DFF_1369_Q_reg ( .D(g30361), .SI(g2661), .SE(test_se), .CLK(CK), .Q(
        g1988), .QN(n5783) );
  SDFFX1 DFF_1370_Q_reg ( .D(g25705), .SI(g1988), .SE(test_se), .CLK(CK), .Q(
        test_so96), .QN(n5427) );
  SDFFX1 DFF_1371_Q_reg ( .D(g24260), .SI(test_si97), .SE(test_se), .CLK(CK), 
        .Q(g1548), .QN(n5546) );
  SDFFX1 DFF_1372_Q_reg ( .D(g29257), .SI(g1548), .SE(test_se), .CLK(CK), .Q(
        g3106), .QN(n5742) );
  SDFFX1 DFF_1373_Q_reg ( .D(g34461), .SI(g3106), .SE(test_se), .CLK(CK), .Q(
        g4659), .QN() );
  SDFFX1 DFF_1374_Q_reg ( .D(g34258), .SI(g4659), .SE(test_se), .CLK(CK), .Q(
        g4358), .QN(n5348) );
  SDFFX1 DFF_1375_Q_reg ( .D(g32993), .SI(g4358), .SE(test_se), .CLK(CK), .Q(
        g1792), .QN(n5359) );
  SDFFX1 DFF_1376_Q_reg ( .D(g33992), .SI(g1792), .SE(test_se), .CLK(CK), .Q(
        g2084), .QN() );
  SDFFX1 DFF_1378_Q_reg ( .D(g30394), .SI(g2084), .SE(test_se), .CLK(CK), .Q(
        g3187), .QN() );
  SDFFX1 DFF_1379_Q_reg ( .D(g34449), .SI(g3187), .SE(test_se), .CLK(CK), .Q(
        g4311), .QN(n5323) );
  SDFFX1 DFF_1380_Q_reg ( .D(g34019), .SI(g4311), .SE(test_se), .CLK(CK), .Q(
        g2583), .QN(n5800) );
  SDFFX1 DFF_1381_Q_reg ( .D(g18597), .SI(g2583), .SE(test_se), .CLK(CK), .Q(
        n9240), .QN(DFF_1381_n1) );
  SDFFX1 DFF_1382_Q_reg ( .D(g29231), .SI(n9240), .SE(test_se), .CLK(CK), .Q(
        g1094), .QN(n5697) );
  SDFFX1 DFF_1383_Q_reg ( .D(g25682), .SI(g1094), .SE(test_se), .CLK(CK), .Q(
        test_so97), .QN(n5448) );
  SDFFX1 DFF_1384_Q_reg ( .D(g21897), .SI(test_si98), .SE(test_se), .CLK(CK), 
        .Q(g4284), .QN() );
  SDFFX1 DFF_1386_Q_reg ( .D(g30395), .SI(g4284), .SE(test_se), .CLK(CK), .Q(
        g3191), .QN() );
  SDFFX1 DFF_1387_Q_reg ( .D(g21892), .SI(g3191), .SE(test_se), .CLK(CK), .Q(
        g4239), .QN() );
  SDFFX1 DFF_1389_Q_reg ( .D(g8789), .SI(g4239), .SE(test_se), .CLK(CK), .Q(
        g4180), .QN(n5380) );
  SDFFX1 DFF_1390_Q_reg ( .D(g28048), .SI(g4180), .SE(test_se), .CLK(CK), .Q(
        g691), .QN(n5520) );
  SDFFX1 DFF_1391_Q_reg ( .D(g34723), .SI(g691), .SE(test_se), .CLK(CK), .Q(
        g534), .QN(n5490) );
  SDFFX1 DFF_1393_Q_reg ( .D(g25598), .SI(g534), .SE(test_se), .CLK(CK), .Q(
        g385), .QN(n5632) );
  SDFFX1 DFF_1394_Q_reg ( .D(g33987), .SI(g385), .SE(test_se), .CLK(CK), .Q(
        g2004), .QN(n5818) );
  SDFFX1 DFF_1395_Q_reg ( .D(g30380), .SI(g2004), .SE(test_se), .CLK(CK), .Q(
        g2527), .QN(n5420) );
  SDFFX1 DFF_1396_Q_reg ( .D(g9555), .SI(g2527), .SE(test_se), .CLK(CK), .Q(
        g5456), .QN() );
  SDFFX1 DFF_1397_Q_reg ( .D(g26965), .SI(g5456), .SE(test_se), .CLK(CK), .Q(
        n6007), .QN() );
  SDFFX1 DFF_1398_Q_reg ( .D(g25706), .SI(n6007), .SE(test_se), .CLK(CK), .Q(
        test_so98), .QN(n5444) );
  SDFFX1 DFF_1399_Q_reg ( .D(g30458), .SI(test_si99), .SE(test_se), .CLK(CK), 
        .Q(g4507), .QN(n5846) );
  SDFFX1 DFF_1400_Q_reg ( .D(g24338), .SI(g4507), .SE(test_se), .CLK(CK), .Q(
        g5348), .QN() );
  SDFFX1 DFF_1401_Q_reg ( .D(g30400), .SI(g5348), .SE(test_se), .CLK(CK), .Q(
        g3223), .QN() );
  SDFFX1 DFF_1403_Q_reg ( .D(g34623), .SI(g3223), .SE(test_se), .CLK(CK), .Q(
        g2970), .QN() );
  SDFFX1 DFF_1404_Q_reg ( .D(g24343), .SI(g2970), .SE(test_se), .CLK(CK), .Q(
        g5698), .QN() );
  SDFFX1 DFF_1406_Q_reg ( .D(g30473), .SI(g5698), .SE(test_se), .CLK(CK), .Q(
        g5260), .QN() );
  SDFFX1 DFF_1407_Q_reg ( .D(g24252), .SI(g5260), .SE(test_se), .CLK(CK), .Q(
        g1521), .QN(n5577) );
  SDFFX1 DFF_1408_Q_reg ( .D(g33028), .SI(g1521), .SE(test_se), .CLK(CK), .Q(
        g3522), .QN(n5383) );
  SDFFX1 DFF_1409_Q_reg ( .D(g29258), .SI(g3522), .SE(test_se), .CLK(CK), .Q(
        g3115), .QN() );
  SDFFX1 DFF_1410_Q_reg ( .D(g30407), .SI(g3115), .SE(test_se), .CLK(CK), .Q(
        g3251), .QN() );
  SDFFX1 DFF_1411_Q_reg ( .D(g26958), .SI(g3251), .SE(test_se), .CLK(CK), .Q(
        g12832), .QN() );
  SDFFX1 DFF_1412_Q_reg ( .D(g34457), .SI(g12832), .SE(test_se), .CLK(CK), .Q(
        test_so99), .QN(n5309) );
  SDFFX1 DFF_1413_Q_reg ( .D(g33568), .SI(test_si100), .SE(test_se), .CLK(CK), 
        .Q(g1996), .QN(n5355) );
  SDFFX1 DFF_1414_Q_reg ( .D(g25663), .SI(g1996), .SE(test_se), .CLK(CK), .Q(
        g8342), .QN() );
  SDFFX1 DFF_1415_Q_reg ( .D(g26964), .SI(g8342), .SE(test_se), .CLK(CK), .Q(
        g4515), .QN() );
  SDFFX1 DFF_1416_Q_reg ( .D(g8786), .SI(g4515), .SE(test_se), .CLK(CK), .Q(
        g8787), .QN() );
  SDFFX1 DFF_1417_Q_reg ( .D(g34735), .SI(g8787), .SE(test_se), .CLK(CK), .Q(
        g4300), .QN(n5639) );
  SDFFX1 DFF_1418_Q_reg ( .D(g30352), .SI(g4300), .SE(test_se), .CLK(CK), .Q(
        n9236), .QN(n5626) );
  SDFFX1 DFF_1419_Q_reg ( .D(g33543), .SI(n9236), .SE(test_se), .CLK(CK), .Q(
        g1379), .QN() );
  SDFFX1 DFF_1420_Q_reg ( .D(g24271), .SI(g1379), .SE(test_se), .CLK(CK), .Q(
        g11388), .QN(n5433) );
  SDFFX1 DFF_1422_Q_reg ( .D(g33981), .SI(g11388), .SE(test_se), .CLK(CK), .Q(
        g1878), .QN(n5793) );
  SDFFX1 DFF_1423_Q_reg ( .D(g30500), .SI(g1878), .SE(test_se), .CLK(CK), .Q(
        g5619), .QN() );
  SDFFX1 DFF_1424_Q_reg ( .D(g34649), .SI(g5619), .SE(test_se), .CLK(CK), .Q(
        g71), .QN() );
  SDFFX1 DFF_1425_Q_reg ( .D(g29277), .SI(g71), .SE(test_se), .CLK(CK), .Q(
        g20049), .QN() );
  SDFFX1 DFF_748_Q_reg ( .D(n1461), .SI(g4704), .SE(test_se), .CLK(CK), .Q(g22), .QN() );
  SDFFX1 DFF_591_Q_reg ( .D(g25612), .SI(g3897), .SE(test_se), .CLK(CK), .Q(
        g518), .QN(n5287) );
  SDFFX1 DFF_845_Q_reg ( .D(g28060), .SI(g626), .SE(test_se), .CLK(CK), .Q(
        g2729), .QN() );
  OA22X1 U5132 ( .IN1(n1277), .IN2(1'b1), .IN3(n2502), .IN4(n2455), .Q(n2500)
         );
  OA22X1 U5133 ( .IN1(n1452), .IN2(1'b1), .IN3(n2505), .IN4(n1423), .Q(n2504)
         );
  OA221X1 U5134 ( .IN1(test_so52), .IN2(g939), .IN3(n1309), .IN4(1'b1), .IN5(
        n6211), .Q(n2503) );
  OA221X1 U5135 ( .IN1(g209), .IN2(g538), .IN3(n1457), .IN4(1'b1), .IN5(n6227), 
        .Q(g34719) );
  OA221X1 U5136 ( .IN1(g546), .IN2(n5520), .IN3(n1455), .IN4(1'b1), .IN5(n6233), .Q(n2512) );
  OA221X1 U5137 ( .IN1(g199), .IN2(g222), .IN3(n1277), .IN4(1'b1), .IN5(n6214), 
        .Q(n2513) );
  OA221X1 U5138 ( .IN1(g550), .IN2(n5657), .IN3(n1452), .IN4(1'b1), .IN5(n6216), .Q(n2514) );
  OA221X1 U5139 ( .IN1(g301), .IN2(g534), .IN3(n1453), .IN4(1'b1), .IN5(n6213), 
        .Q(n2510) );
  OA22X1 U5140 ( .IN1(n1277), .IN2(1'b1), .IN3(n2496), .IN4(n2453), .Q(n2494)
         );
  OA22X1 U5141 ( .IN1(n1452), .IN2(1'b1), .IN3(n2499), .IN4(n2447), .Q(n2498)
         );
  OA221X1 U5142 ( .IN1(g1277), .IN2(g1283), .IN3(n1309), .IN4(1'b1), .IN5(
        n6210), .Q(n2497) );
  OA221X1 U5143 ( .IN1(test_so14), .IN2(test_so74), .IN3(1'b1), .IN4(n2461), 
        .IN5(n6222), .Q(n2460) );
  OA221X1 U5144 ( .IN1(g4153), .IN2(g4172), .IN3(n1453), .IN4(1'b1), .IN5(
        n6218), .Q(g34733) );
  OA221X1 U5145 ( .IN1(g4072), .IN2(g4176), .IN3(n1452), .IN4(1'b1), .IN5(
        n6205), .Q(n2490) );
  OA221X1 U5146 ( .IN1(g2932), .IN2(g2999), .IN3(n1456), .IN4(1'b1), .IN5(
        n6224), .Q(g34805) );
  OA221X1 U5147 ( .IN1(g2890), .IN2(n5928), .IN3(n1277), .IN4(1'b1), .IN5(
        n6226), .Q(n2462) );
  OA221X1 U5148 ( .IN1(test_so63), .IN2(g4300), .IN3(n1453), .IN4(1'b1), .IN5(
        n6206), .Q(n2488) );
  OA221X1 U5149 ( .IN1(g2864), .IN2(n2437), .IN3(n1455), .IN4(1'b1), .IN5(
        n6208), .Q(n2472) );
  OA221X1 U5150 ( .IN1(g2898), .IN2(n2438), .IN3(n1454), .IN4(1'b1), .IN5(
        n6219), .Q(n2468) );
  OA221X1 U5151 ( .IN1(g2886), .IN2(g2946), .IN3(n1309), .IN4(1'b1), .IN5(
        n6212), .Q(n2463) );
  OA221X1 U5152 ( .IN1(n2441), .IN2(n2483), .IN3(n1457), .IN4(1'b1), .IN5(
        n6207), .Q(n2482) );
  OA221X1 U5153 ( .IN1(g2878), .IN2(n5926), .IN3(n1452), .IN4(1'b1), .IN5(
        n6598), .Q(n2465) );
  OA221X1 U5154 ( .IN1(n2432), .IN2(n2467), .IN3(n1453), .IN4(1'b1), .IN5(
        n6209), .Q(n2466) );
  OA221X1 U5155 ( .IN1(n2439), .IN2(n2481), .IN3(n1456), .IN4(1'b1), .IN5(
        n6215), .Q(n2480) );
  OA221X1 U5156 ( .IN1(n5928), .IN2(n2451), .IN3(n1455), .IN4(1'b1), .IN5(
        n6223), .Q(n2450) );
  OA221X1 U5157 ( .IN1(n1453), .IN2(1'b1), .IN3(n2435), .IN4(n2436), .IN5(
        n6225), .Q(n2434) );
  OA221X1 U5158 ( .IN1(g2941), .IN2(n2444), .IN3(n1454), .IN4(1'b1), .IN5(
        n6230), .Q(n2443) );
  OA221X1 U5159 ( .IN1(n2447), .IN2(n2448), .IN3(n1309), .IN4(1'b1), .IN5(
        n6220), .Q(n2446) );
  OA221X1 U5160 ( .IN1(n2457), .IN2(n2458), .IN3(n1457), .IN4(1'b1), .IN5(
        n6217), .Q(n2456) );
  OA221X1 U5161 ( .IN1(n2453), .IN2(n2454), .IN3(n1456), .IN4(1'b1), .IN5(
        n6234), .Q(n2452) );
  AO221X1 U5162 ( .IN1(n2396), .IN2(1'b0), .IN3(n5842), .IN4(n2397), .IN5(
        n6084), .Q(n2395) );
  AO22X1 U5163 ( .IN1(n2540), .IN2(1'b0), .IN3(n2551), .IN4(n6289), .Q(g34601)
         );
  NOR2X0 U5164 ( .IN1(1'b0), .IN2(n5286), .QN(n2551) );
  NOR2X0 U5165 ( .IN1(n6082), .IN2(1'b0), .QN(n2538) );
  AO222X1 U5166 ( .IN1(n2538), .IN2(g2950), .IN3(n2540), .IN4(1'b0), .IN5(
        g2936), .IN6(n6105), .Q(g34621) );
  AO222X1 U5167 ( .IN1(n2538), .IN2(test_so1), .IN3(1'b0), .IN4(n2521), .IN5(
        g2984), .IN6(n6104), .Q(g34617) );
  AO222X1 U5168 ( .IN1(n2538), .IN2(test_so22), .IN3(1'b0), .IN4(n2535), .IN5(
        g2950), .IN6(n6105), .Q(g34622) );
  AO222X1 U5169 ( .IN1(1'b0), .IN2(n2518), .IN3(n2538), .IN4(g2936), .IN5(
        g2922), .IN6(n6104), .Q(g34620) );
  AO222X1 U5170 ( .IN1(n2538), .IN2(g2922), .IN3(1'b0), .IN4(n2523), .IN5(
        g2912), .IN6(n6104), .Q(g34619) );
  AO222X1 U5171 ( .IN1(n2538), .IN2(g2912), .IN3(1'b0), .IN4(n2522), .IN5(
        test_so1), .IN6(n6104), .Q(g34618) );
  AO222X1 U5172 ( .IN1(n2538), .IN2(g2970), .IN3(1'b0), .IN4(n2534), .IN5(
        test_so22), .IN6(n6089), .Q(g34623) );
  MUX21X2 U5173 ( .IN1(n2544), .IN2(test_so95), .S(n6102), .Q(g34613) );
  NOR2X0 U5174 ( .IN1(g23002), .IN2(1'b0), .QN(n2544) );
  MUX21X2 U5175 ( .IN1(n2543), .IN2(g37), .S(n6103), .Q(g34614) );
  NOR2X0 U5176 ( .IN1(1'b0), .IN2(n5342), .QN(n2543) );
  AO22X1 U5177 ( .IN1(n2516), .IN2(test_so45), .IN3(n2522), .IN4(1'b0), .Q(
        g34626) );
  NOR2X0 U5178 ( .IN1(n6081), .IN2(1'b0), .QN(n2516) );
  AO22X1 U5179 ( .IN1(n2516), .IN2(g3853), .IN3(n2521), .IN4(1'b0), .Q(g34627)
         );
  AO22X1 U5180 ( .IN1(n2516), .IN2(g3151), .IN3(n2523), .IN4(1'b0), .Q(g34625)
         );
  AO22X1 U5181 ( .IN1(n2516), .IN2(g6545), .IN3(1'b0), .IN4(n2518), .Q(g34647)
         );
  AO22X1 U5182 ( .IN1(n2516), .IN2(g2689), .IN3(n2535), .IN4(1'b0), .Q(g34606)
         );
  AO222X1 U5183 ( .IN1(n2516), .IN2(g2704), .IN3(n2532), .IN4(1'b0), .IN5(
        g2697), .IN6(n6099), .Q(g34608) );
  AO222X1 U5184 ( .IN1(n2516), .IN2(g2697), .IN3(n2534), .IN4(1'b0), .IN5(
        g2689), .IN6(n6099), .Q(g34607) );
  AO22X1 U5185 ( .IN1(n2519), .IN2(g5853), .IN3(n2522), .IN4(1'b0), .Q(g34645)
         );
  NOR2X0 U5186 ( .IN1(n6080), .IN2(1'b0), .QN(n2519) );
  AO22X1 U5187 ( .IN1(1'b0), .IN2(n2518), .IN3(n2519), .IN4(g5160), .Q(g34643)
         );
  AO22X1 U5188 ( .IN1(n2519), .IN2(g6199), .IN3(1'b0), .IN4(n2521), .Q(g34646)
         );
  AO22X1 U5189 ( .IN1(n2519), .IN2(g5507), .IN3(n2523), .IN4(1'b0), .Q(g34644)
         );
  AO22X1 U5190 ( .IN1(n2519), .IN2(g2130), .IN3(n2535), .IN4(1'b0), .Q(g34603)
         );
  AO222X1 U5191 ( .IN1(n2519), .IN2(g2145), .IN3(n2532), .IN4(1'b0), .IN5(
        g2138), .IN6(n6098), .Q(g34605) );
  AO222X1 U5192 ( .IN1(n2519), .IN2(g2138), .IN3(n2534), .IN4(1'b0), .IN5(
        g2130), .IN6(n6098), .Q(g34604) );
  NOR2X0 U5193 ( .IN1(n6082), .IN2(1'b0), .QN(n2537) );
  AO222X1 U5194 ( .IN1(n2521), .IN2(1'b0), .IN3(n2537), .IN4(g2844), .IN5(
        g2890), .IN6(n6099), .Q(g34609) );
  AO222X1 U5195 ( .IN1(n2522), .IN2(1'b0), .IN3(n2537), .IN4(g2852), .IN5(
        g2844), .IN6(n6100), .Q(g34610) );
  AO222X1 U5196 ( .IN1(n2523), .IN2(1'b0), .IN3(n2537), .IN4(g2860), .IN5(
        g2852), .IN6(n6100), .Q(g34611) );
  AO222X1 U5197 ( .IN1(n2518), .IN2(1'b0), .IN3(n2537), .IN4(test_so95), .IN5(
        g2860), .IN6(n6102), .Q(g34612) );
  AO222X1 U5198 ( .IN1(n2537), .IN2(g4157), .IN3(n2532), .IN4(1'b0), .IN5(
        g4146), .IN6(n6090), .Q(g34629) );
  AO222X1 U5199 ( .IN1(n2537), .IN2(g4146), .IN3(n2534), .IN4(1'b0), .IN5(
        g4176), .IN6(n6090), .Q(g34628) );
  NOR2X0 U5200 ( .IN1(n6083), .IN2(1'b0), .QN(n2492) );
  AO222X1 U5201 ( .IN1(n2535), .IN2(1'b0), .IN3(n2492), .IN4(g2873), .IN5(
        g2868), .IN6(n6104), .Q(g34615) );
  AO222X1 U5202 ( .IN1(g2994), .IN2(n2492), .IN3(n2493), .IN4(1'b0), .IN5(
        g2999), .IN6(n6095), .Q(g34732) );
  AO222X1 U5203 ( .IN1(n2492), .IN2(g2868), .IN3(n2540), .IN4(1'b0), .IN5(
        g2988), .IN6(n6104), .Q(g34616) );
  AO222X1 U5204 ( .IN1(n2518), .IN2(1'b0), .IN3(n2492), .IN4(g2988), .IN5(
        g2994), .IN6(n6089), .Q(g34624) );
  NOR2X0 U5205 ( .IN1(n6083), .IN2(1'b0), .QN(n2529) );
  AO22X1 U5206 ( .IN1(1'b0), .IN2(n2521), .IN3(n2529), .IN4(g4727), .Q(g34633)
         );
  AO222X1 U5207 ( .IN1(1'b0), .IN2(n2518), .IN3(n2529), .IN4(g4722), .IN5(
        g4717), .IN6(n6092), .Q(g34636) );
  AO222X1 U5208 ( .IN1(1'b0), .IN2(n2522), .IN3(n2529), .IN4(g4732), .IN5(
        g4727), .IN6(n6092), .Q(g34634) );
  AO222X1 U5209 ( .IN1(1'b0), .IN2(n2523), .IN3(n2529), .IN4(g4717), .IN5(
        g4732), .IN6(n6092), .Q(g34635) );
  AO222X1 U5210 ( .IN1(g4737), .IN2(n2529), .IN3(n2525), .IN4(1'b0), .IN5(
        g4722), .IN6(n6092), .Q(g34637) );
  NOR2X0 U5211 ( .IN1(n6083), .IN2(1'b0), .QN(n2533) );
  AO222X1 U5212 ( .IN1(n2535), .IN2(1'b0), .IN3(n2533), .IN4(g4253), .IN5(
        g4300), .IN6(n6091), .Q(g34630) );
  AO222X1 U5213 ( .IN1(n2534), .IN2(1'b0), .IN3(n2533), .IN4(test_so67), .IN5(
        g4253), .IN6(n6091), .Q(g34631) );
  AO222X1 U5214 ( .IN1(n2532), .IN2(1'b0), .IN3(n2533), .IN4(g4245), .IN5(
        test_so67), .IN6(n6091), .Q(g34632) );
  NOR2X0 U5215 ( .IN1(n6083), .IN2(1'b0), .QN(n2524) );
  AO22X1 U5216 ( .IN1(1'b0), .IN2(n2521), .IN3(n2524), .IN4(g4917), .Q(g34638)
         );
  AO222X1 U5217 ( .IN1(1'b0), .IN2(n2518), .IN3(n2524), .IN4(g4912), .IN5(
        g4907), .IN6(n6094), .Q(g34641) );
  AO222X1 U5218 ( .IN1(1'b0), .IN2(n2522), .IN3(n2524), .IN4(g4922), .IN5(
        g4917), .IN6(n6093), .Q(g34639) );
  AO222X1 U5219 ( .IN1(1'b0), .IN2(n2523), .IN3(n2524), .IN4(g4907), .IN5(
        g4922), .IN6(n6094), .Q(g34640) );
  AO222X1 U5220 ( .IN1(g4927), .IN2(n2524), .IN3(n2525), .IN4(1'b0), .IN5(
        g4912), .IN6(n6094), .Q(g34642) );
  AO21X1 U5221 ( .IN1(n3177), .IN2(n2172), .IN3(g24183), .Q(n2884) );
  AOI21X1 U5222 ( .IN1(n3254), .IN2(n2172), .IN3(g24183), .QN(n2978) );
  AO21X1 U5223 ( .IN1(g24169), .IN2(n5634), .IN3(n2416), .Q(n2414) );
  AND2X1 U5224 ( .IN1(g24174), .IN2(n2668), .Q(n2714) );
  AO21X1 U5225 ( .IN1(g24172), .IN2(g37), .IN3(g24183), .Q(n2668) );
  AND3X1 U5226 ( .IN1(g24168), .IN2(n5605), .IN3(n4670), .Q(n3719) );
  INVX0 U5227 ( .IN(n4169), .QN(n1548) );
  INVX0 U5228 ( .IN(n4187), .QN(n1583) );
  AO221X1 U5229 ( .IN1(g2453), .IN2(n1392), .IN3(g2461), .IN4(n6086), .IN5(
        n3540), .Q(g33011) );
  AO22X1 U5230 ( .IN1(g3451), .IN2(n6125), .IN3(n5038), .IN4(n6297), .Q(g25664) );
  AO221X1 U5231 ( .IN1(g2028), .IN2(n1395), .IN3(test_so59), .IN4(n6085), 
        .IN5(n3597), .Q(g32999) );
  AO221X1 U5232 ( .IN1(g1624), .IN2(n1398), .IN3(g1632), .IN4(n6085), .IN5(
        n3650), .Q(g32987) );
  AO221X1 U5233 ( .IN1(g2185), .IN2(n1394), .IN3(g2193), .IN4(n6085), .IN5(
        n3578), .Q(g33003) );
  AO22X1 U5234 ( .IN1(g6148), .IN2(n6124), .IN3(n4995), .IN4(n6299), .Q(g25744) );
  AO22X1 U5235 ( .IN1(g6494), .IN2(n6124), .IN3(n4990), .IN4(n6298), .Q(g25758) );
  AO221X1 U5236 ( .IN1(g1894), .IN2(n1396), .IN3(g1902), .IN4(n6087), .IN5(
        n3615), .Q(g32995) );
  AO221X1 U5237 ( .IN1(g2587), .IN2(n1391), .IN3(test_so34), .IN4(n6086), 
        .IN5(n3521), .Q(g33015) );
  AO221X1 U5238 ( .IN1(g1760), .IN2(n1397), .IN3(g1768), .IN4(n6084), .IN5(
        n3632), .Q(g32991) );
  AO22X1 U5239 ( .IN1(g5456), .IN2(n6124), .IN3(n5005), .IN4(n6299), .Q(g25716) );
  AO22X1 U5240 ( .IN1(g3802), .IN2(n6125), .IN3(n5033), .IN4(n6298), .Q(g25678) );
  AO22X1 U5241 ( .IN1(g5802), .IN2(n6124), .IN3(n5000), .IN4(n6295), .Q(g25730) );
  AO221X1 U5242 ( .IN1(g2319), .IN2(n1393), .IN3(g2327), .IN4(n6085), .IN5(
        n3559), .Q(g33007) );
  AO22X1 U5243 ( .IN1(g3100), .IN2(n6126), .IN3(n5043), .IN4(n6293), .Q(g25650) );
  AO22X1 U5244 ( .IN1(g20901), .IN2(n6122), .IN3(n2983), .IN4(n6280), .Q(
        g33963) );
  AO22X1 U5245 ( .IN1(n6135), .IN2(g4122), .IN3(n3935), .IN4(n6281), .Q(g30457) );
  INVX0 U5246 ( .IN(g6753), .QN(n5894) );
  INVX0 U5247 ( .IN(n5894), .QN(g18092) );
  INVX0 U5248 ( .IN(g6751), .QN(n5896) );
  INVX0 U5249 ( .IN(n5896), .QN(g18100) );
  INVX0 U5250 ( .IN(g6747), .QN(n5898) );
  INVX0 U5251 ( .IN(n5898), .QN(g18097) );
  INVX0 U5252 ( .IN(g6746), .QN(n5900) );
  INVX0 U5253 ( .IN(n5900), .QN(g18101) );
  INVX0 U5254 ( .IN(g36), .QN(n5902) );
  INVX0 U5255 ( .IN(n5902), .QN(g21698) );
  INVX0 U5256 ( .IN(g6745), .QN(n5904) );
  INVX0 U5257 ( .IN(n5904), .QN(g18099) );
  INVX0 U5258 ( .IN(g64), .QN(n5906) );
  INVX0 U5259 ( .IN(n5906), .QN(g24165) );
  INVX0 U5260 ( .IN(g125), .QN(n5908) );
  INVX0 U5261 ( .IN(n5908), .QN(g24180) );
  INVX0 U5262 ( .IN(g120), .QN(n5910) );
  INVX0 U5263 ( .IN(n5910), .QN(g24178) );
  INVX0 U5264 ( .IN(g114), .QN(n5912) );
  INVX0 U5265 ( .IN(n5912), .QN(g24175) );
  INVX0 U5266 ( .IN(g6744), .QN(n5914) );
  INVX0 U5267 ( .IN(n5914), .QN(g18098) );
  INVX0 U5268 ( .IN(g124), .QN(n5916) );
  INVX0 U5269 ( .IN(n5916), .QN(g24179) );
  INVX0 U5270 ( .IN(g116), .QN(n5918) );
  INVX0 U5271 ( .IN(n5918), .QN(g24177) );
  INVX0 U5272 ( .IN(g100), .QN(n5920) );
  INVX0 U5273 ( .IN(n5920), .QN(g24173) );
  INVX0 U5274 ( .IN(g99), .QN(n5922) );
  INVX0 U5275 ( .IN(n5922), .QN(g24172) );
  INVX0 U5276 ( .IN(g90), .QN(n5924) );
  INVX0 U5277 ( .IN(n5924), .QN(g24169) );
  INVX0 U5278 ( .IN(g91), .QN(n5926) );
  INVX0 U5279 ( .IN(n5926), .QN(g24170) );
  INVX0 U5280 ( .IN(g44), .QN(n5928) );
  INVX0 U5281 ( .IN(n5928), .QN(g24185) );
  INVX0 U5282 ( .IN(g57), .QN(n5930) );
  INVX0 U5283 ( .IN(n5930), .QN(g24164) );
  INVX0 U5284 ( .IN(g135), .QN(n5932) );
  INVX0 U5285 ( .IN(n5932), .QN(g24184) );
  INVX0 U5286 ( .IN(g92), .QN(n5934) );
  INVX0 U5287 ( .IN(n5934), .QN(g24171) );
  INVX0 U5288 ( .IN(g127), .QN(n5936) );
  INVX0 U5289 ( .IN(n5936), .QN(g24182) );
  INVX0 U5290 ( .IN(g126), .QN(n5938) );
  INVX0 U5291 ( .IN(n5938), .QN(g24181) );
  INVX0 U5292 ( .IN(g115), .QN(n5940) );
  INVX0 U5293 ( .IN(n5940), .QN(g24176) );
  INVX0 U5294 ( .IN(g6750), .QN(n5942) );
  INVX0 U5295 ( .IN(n5942), .QN(g18096) );
  INVX0 U5296 ( .IN(g6749), .QN(n5944) );
  INVX0 U5297 ( .IN(n5944), .QN(g18095) );
  INVX0 U5298 ( .IN(g6748), .QN(n5946) );
  INVX0 U5299 ( .IN(n5946), .QN(g18094) );
  INVX0 U5300 ( .IN(g53), .QN(n5948) );
  INVX0 U5301 ( .IN(n5948), .QN(g24161) );
  INVX0 U5302 ( .IN(g84), .QN(n5950) );
  INVX0 U5303 ( .IN(n5950), .QN(g24168) );
  INVX0 U5304 ( .IN(g134), .QN(n5952) );
  INVX0 U5305 ( .IN(n5952), .QN(g24183) );
  INVX0 U5306 ( .IN(g54), .QN(n5954) );
  INVX0 U5307 ( .IN(n5954), .QN(g24162) );
  INVX0 U5308 ( .IN(g56), .QN(n5956) );
  INVX0 U5309 ( .IN(n5956), .QN(g24163) );
  INVX0 U5310 ( .IN(g113), .QN(n5958) );
  INVX0 U5311 ( .IN(n5958), .QN(g24174) );
  INVX0 U5312 ( .IN(n6580), .QN(n6498) );
  INVX0 U5313 ( .IN(n6660), .QN(n6639) );
  INVX0 U5314 ( .IN(n2930), .QN(n1365) );
  INVX0 U5315 ( .IN(n2953), .QN(n1356) );
  INVX0 U5316 ( .IN(n2906), .QN(n1374) );
  INVX0 U5317 ( .IN(n2966), .QN(n1347) );
  NAND2X0 U5318 ( .IN1(n6236), .IN2(n3127), .QN(n3129) );
  NAND2X0 U5319 ( .IN1(n6227), .IN2(n3167), .QN(n3169) );
  NAND2X0 U5320 ( .IN1(n6223), .IN2(n3148), .QN(n3150) );
  NAND2X0 U5321 ( .IN1(n6237), .IN2(n3107), .QN(n3109) );
  NAND2X0 U5322 ( .IN1(n6216), .IN2(n3208), .QN(n3210) );
  NAND2X0 U5323 ( .IN1(n6225), .IN2(n3228), .QN(n3230) );
  NAND2X0 U5324 ( .IN1(n6665), .IN2(n3188), .QN(n3190) );
  NAND2X0 U5325 ( .IN1(n6226), .IN2(n3246), .QN(n3248) );
  NAND2X0 U5326 ( .IN1(n2102), .IN2(n1558), .QN(n2688) );
  NAND2X0 U5327 ( .IN1(n2134), .IN2(n1704), .QN(n2667) );
  NAND2X0 U5328 ( .IN1(n2455), .IN2(n2453), .QN(g28041) );
  INVX0 U5329 ( .IN(n6679), .QN(n6674) );
  INVX0 U5330 ( .IN(n3094), .QN(n1489) );
  NOR2X0 U5331 ( .IN1(n2868), .IN2(n3160), .QN(n2870) );
  NOR2X0 U5332 ( .IN1(n2845), .IN2(n3141), .QN(n2847) );
  NOR2X0 U5333 ( .IN1(n2822), .IN2(n3122), .QN(n2824) );
  NOR2X0 U5334 ( .IN1(n2798), .IN2(n3102), .QN(n2800) );
  NOR2X0 U5335 ( .IN1(n5503), .IN2(n1365), .QN(n2923) );
  NOR2X0 U5336 ( .IN1(n5505), .IN2(n1374), .QN(n2899) );
  NOR2X0 U5337 ( .IN1(n5504), .IN2(n1356), .QN(n2946) );
  INVX0 U5338 ( .IN(n4314), .QN(n1558) );
  INVX0 U5339 ( .IN(n4292), .QN(n1704) );
  INVX0 U5340 ( .IN(n2962), .QN(n1351) );
  INVX0 U5341 ( .IN(n2939), .QN(n1360) );
  INVX0 U5342 ( .IN(n2916), .QN(n1369) );
  INVX0 U5343 ( .IN(n2892), .QN(n1378) );
  INVX0 U5344 ( .IN(n2884), .QN(n1342) );
  INVX0 U5345 ( .IN(g72), .QN(n5962) );
  NAND2X0 U5346 ( .IN1(g4785), .IN2(g4709), .QN(n4326) );
  NAND2X0 U5347 ( .IN1(g4975), .IN2(g4899), .QN(n4304) );
  NAND2X0 U5348 ( .IN1(g4688), .IN2(n3012), .QN(n2690) );
  NAND2X0 U5349 ( .IN1(g4878), .IN2(n3013), .QN(n2670) );
  INVX0 U5350 ( .IN(g35), .QN(n6683) );
  LSDNX1 U5351 ( .D(g73), .Q(g24167) );
  LSDNX1 U5352 ( .D(g72), .Q(n6018) );
  ISOLANDX1 U5353 ( .D(n5960), .ISO(n1705), .Q(n4689) );
  AO221X1 U5354 ( .IN1(n2123), .IN2(g6736), .IN3(n2122), .IN4(g6732), .IN5(
        n4691), .Q(n5960) );
  ISOLANDX1 U5355 ( .D(n5961), .ISO(n1560), .Q(n4708) );
  AO221X1 U5356 ( .IN1(g31860), .IN2(g5352), .IN3(n1893), .IN4(g5348), .IN5(
        n4710), .Q(n5961) );
  NAND2X1 U5357 ( .IN1(n5467), .IN2(n5321), .QN(n4837) );
  NAND2X1 U5358 ( .IN1(n5322), .IN2(n5466), .QN(n4836) );
  NAND2X1 U5359 ( .IN1(n3010), .IN2(n3011), .QN(g34783) );
  AND2X1 U5360 ( .IN1(n6261), .IN2(n5963), .Q(n2787) );
  INVX0 U5361 ( .IN(n6261), .QN(n6083) );
  INVX0 U5362 ( .IN(n6237), .QN(n6144) );
  INVX0 U5363 ( .IN(n6261), .QN(n6082) );
  INVX0 U5364 ( .IN(n6266), .QN(n6069) );
  INVX0 U5365 ( .IN(n6260), .QN(n6068) );
  INVX0 U5366 ( .IN(n6262), .QN(n6080) );
  INVX0 U5367 ( .IN(n6241), .QN(n6140) );
  INVX0 U5368 ( .IN(n6240), .QN(n6141) );
  INVX0 U5369 ( .IN(n6238), .QN(n6143) );
  INVX0 U5370 ( .IN(n6239), .QN(n6142) );
  INVX0 U5371 ( .IN(n6236), .QN(n6145) );
  INVX0 U5372 ( .IN(n6260), .QN(n6084) );
  INVX0 U5373 ( .IN(n6259), .QN(n6087) );
  INVX0 U5374 ( .IN(n6259), .QN(n6086) );
  INVX0 U5375 ( .IN(n6260), .QN(n6085) );
  INVX0 U5376 ( .IN(n6259), .QN(n6088) );
  INVX0 U5377 ( .IN(n6251), .QN(n6109) );
  INVX0 U5378 ( .IN(n6253), .QN(n6103) );
  INVX0 U5379 ( .IN(n6251), .QN(n6110) );
  INVX0 U5380 ( .IN(n6256), .QN(n6094) );
  INVX0 U5381 ( .IN(n6252), .QN(n6108) );
  INVX0 U5382 ( .IN(n6251), .QN(n6111) );
  INVX0 U5383 ( .IN(n6252), .QN(n6106) );
  INVX0 U5384 ( .IN(n6254), .QN(n6101) );
  INVX0 U5385 ( .IN(n6253), .QN(n6105) );
  INVX0 U5386 ( .IN(n6255), .QN(n6097) );
  INVX0 U5387 ( .IN(n6254), .QN(n6100) );
  INVX0 U5388 ( .IN(n6255), .QN(n6099) );
  INVX0 U5389 ( .IN(n6256), .QN(n6095) );
  INVX0 U5390 ( .IN(n6252), .QN(n6107) );
  INVX0 U5391 ( .IN(n6257), .QN(n6093) );
  INVX0 U5392 ( .IN(n6254), .QN(n6102) );
  INVX0 U5393 ( .IN(n6250), .QN(n6112) );
  INVX0 U5394 ( .IN(n6255), .QN(n6098) );
  INVX0 U5395 ( .IN(n6258), .QN(n6091) );
  INVX0 U5396 ( .IN(n6253), .QN(n6104) );
  INVX0 U5397 ( .IN(n6256), .QN(n6096) );
  INVX0 U5398 ( .IN(n6250), .QN(n6113) );
  INVX0 U5399 ( .IN(n6250), .QN(n6114) );
  INVX0 U5400 ( .IN(n6257), .QN(n6092) );
  INVX0 U5401 ( .IN(n6258), .QN(n6090) );
  INVX0 U5402 ( .IN(n6258), .QN(n6089) );
  INVX0 U5403 ( .IN(n6249), .QN(n6115) );
  INVX0 U5404 ( .IN(n6249), .QN(n6116) );
  INVX0 U5405 ( .IN(n6262), .QN(n6081) );
  INVX0 U5406 ( .IN(n6249), .QN(n6117) );
  INVX0 U5407 ( .IN(n6248), .QN(n6118) );
  INVX0 U5408 ( .IN(n6264), .QN(n6076) );
  INVX0 U5409 ( .IN(n6266), .QN(n6071) );
  INVX0 U5410 ( .IN(n6267), .QN(n6065) );
  INVX0 U5411 ( .IN(n6262), .QN(n6066) );
  INVX0 U5412 ( .IN(n6263), .QN(n6077) );
  INVX0 U5413 ( .IN(n6263), .QN(n6072) );
  INVX0 U5414 ( .IN(n6265), .QN(n6070) );
  INVX0 U5415 ( .IN(n6264), .QN(n6075) );
  INVX0 U5416 ( .IN(n6267), .QN(n6067) );
  INVX0 U5417 ( .IN(n6266), .QN(n6073) );
  INVX0 U5418 ( .IN(n6265), .QN(n6074) );
  INVX0 U5419 ( .IN(n6263), .QN(n6078) );
  INVX0 U5420 ( .IN(n6265), .QN(n6064) );
  INVX0 U5421 ( .IN(n6264), .QN(n6063) );
  INVX0 U5422 ( .IN(n6248), .QN(n6119) );
  INVX0 U5423 ( .IN(n6248), .QN(n6120) );
  INVX0 U5424 ( .IN(n6247), .QN(n6121) );
  INVX0 U5425 ( .IN(n6257), .QN(n6122) );
  INVX0 U5426 ( .IN(n6261), .QN(n6079) );
  INVX0 U5427 ( .IN(n6245), .QN(n6129) );
  INVX0 U5428 ( .IN(n6247), .QN(n6123) );
  INVX0 U5429 ( .IN(n6245), .QN(n6130) );
  INVX0 U5430 ( .IN(n6246), .QN(n6127) );
  INVX0 U5431 ( .IN(n6244), .QN(n6132) );
  INVX0 U5432 ( .IN(n6246), .QN(n6126) );
  INVX0 U5433 ( .IN(n6244), .QN(n6133) );
  INVX0 U5434 ( .IN(n6246), .QN(n6125) );
  INVX0 U5435 ( .IN(n6244), .QN(n6131) );
  INVX0 U5436 ( .IN(n6247), .QN(n6124) );
  INVX0 U5437 ( .IN(n6245), .QN(n6128) );
  INVX0 U5438 ( .IN(n6243), .QN(n6134) );
  INVX0 U5439 ( .IN(n6243), .QN(n6135) );
  INVX0 U5440 ( .IN(n6243), .QN(n6136) );
  INVX0 U5441 ( .IN(n6242), .QN(n6137) );
  INVX0 U5442 ( .IN(n6242), .QN(n6138) );
  INVX0 U5443 ( .IN(n6242), .QN(n6139) );
  INVX0 U5444 ( .IN(n6235), .QN(n6146) );
  INVX0 U5445 ( .IN(n6498), .QN(n6261) );
  INVX0 U5446 ( .IN(n6510), .QN(n6237) );
  INVX0 U5447 ( .IN(n6495), .QN(n6266) );
  INVX0 U5448 ( .IN(n6497), .QN(n6262) );
  INVX0 U5449 ( .IN(n6498), .QN(n6260) );
  INVX0 U5450 ( .IN(n6452), .QN(n6353) );
  INVX0 U5451 ( .IN(n6450), .QN(n6357) );
  INVX0 U5452 ( .IN(n6448), .QN(n6360) );
  INVX0 U5453 ( .IN(n6442), .QN(n6372) );
  INVX0 U5454 ( .IN(n6520), .QN(n6211) );
  INVX0 U5455 ( .IN(n6519), .QN(n6214) );
  INVX0 U5456 ( .IN(n6517), .QN(n6218) );
  INVX0 U5457 ( .IN(n6511), .QN(n6233) );
  INVX0 U5458 ( .IN(n6519), .QN(n6213) );
  INVX0 U5459 ( .IN(n6513), .QN(n6227) );
  INVX0 U5460 ( .IN(n6518), .QN(n6216) );
  INVX0 U5461 ( .IN(n6628), .QN(n6229) );
  INVX0 U5462 ( .IN(n6513), .QN(n6228) );
  INVX0 U5463 ( .IN(n6512), .QN(n6230) );
  INVX0 U5464 ( .IN(n6517), .QN(n6217) );
  INVX0 U5465 ( .IN(n6528), .QN(n6220) );
  INVX0 U5466 ( .IN(n6511), .QN(n6232) );
  INVX0 U5467 ( .IN(n6453), .QN(n6219) );
  INVX0 U5468 ( .IN(n6515), .QN(n6223) );
  INVX0 U5469 ( .IN(n6514), .QN(n6226) );
  INVX0 U5470 ( .IN(n6516), .QN(n6222) );
  INVX0 U5471 ( .IN(n6629), .QN(n6234) );
  INVX0 U5472 ( .IN(n6518), .QN(n6215) );
  INVX0 U5473 ( .IN(n6516), .QN(n6221) );
  INVX0 U5474 ( .IN(n6520), .QN(n6212) );
  INVX0 U5475 ( .IN(n6514), .QN(n6225) );
  INVX0 U5476 ( .IN(n6512), .QN(n6231) );
  INVX0 U5477 ( .IN(n6515), .QN(n6224) );
  INVX0 U5478 ( .IN(n6510), .QN(n6236) );
  INVX0 U5479 ( .IN(n6624), .QN(n6235) );
  INVX0 U5480 ( .IN(n6509), .QN(n6238) );
  INVX0 U5481 ( .IN(n6508), .QN(n6240) );
  INVX0 U5482 ( .IN(n6508), .QN(n6241) );
  INVX0 U5483 ( .IN(n6509), .QN(n6239) );
  INVX0 U5484 ( .IN(n6496), .QN(n6264) );
  INVX0 U5485 ( .IN(n6504), .QN(n6248) );
  INVX0 U5486 ( .IN(n6496), .QN(n6265) );
  INVX0 U5487 ( .IN(n6497), .QN(n6263) );
  INVX0 U5488 ( .IN(n6504), .QN(n6249) );
  INVX0 U5489 ( .IN(n6507), .QN(n6242) );
  INVX0 U5490 ( .IN(n6503), .QN(n6251) );
  INVX0 U5491 ( .IN(n6499), .QN(n6259) );
  INVX0 U5492 ( .IN(n6505), .QN(n6246) );
  INVX0 U5493 ( .IN(n6502), .QN(n6252) );
  INVX0 U5494 ( .IN(n6506), .QN(n6244) );
  INVX0 U5495 ( .IN(n6507), .QN(n6243) );
  INVX0 U5496 ( .IN(n6501), .QN(n6254) );
  INVX0 U5497 ( .IN(n6505), .QN(n6247) );
  INVX0 U5498 ( .IN(n6501), .QN(n6255) );
  INVX0 U5499 ( .IN(n6502), .QN(n6253) );
  INVX0 U5500 ( .IN(n6500), .QN(n6256) );
  INVX0 U5501 ( .IN(n6503), .QN(n6250) );
  INVX0 U5502 ( .IN(n6506), .QN(n6245) );
  INVX0 U5503 ( .IN(n6500), .QN(n6257) );
  INVX0 U5504 ( .IN(n6499), .QN(n6258) );
  INVX0 U5505 ( .IN(n6495), .QN(n6267) );
  INVX0 U5506 ( .IN(n6494), .QN(n6269) );
  INVX0 U5507 ( .IN(n6492), .QN(n6273) );
  INVX0 U5508 ( .IN(n6493), .QN(n6270) );
  INVX0 U5509 ( .IN(n6494), .QN(n6268) );
  INVX0 U5510 ( .IN(n6492), .QN(n6272) );
  INVX0 U5511 ( .IN(n6493), .QN(n6271) );
  INVX0 U5512 ( .IN(n6491), .QN(n6274) );
  INVX0 U5513 ( .IN(n6491), .QN(n6275) );
  INVX0 U5514 ( .IN(n6490), .QN(n6276) );
  INVX0 U5515 ( .IN(n6484), .QN(n6288) );
  INVX0 U5516 ( .IN(n6485), .QN(n6287) );
  INVX0 U5517 ( .IN(n6483), .QN(n6290) );
  INVX0 U5518 ( .IN(n6489), .QN(n6279) );
  INVX0 U5519 ( .IN(n6484), .QN(n6289) );
  INVX0 U5520 ( .IN(n6481), .QN(n6295) );
  INVX0 U5521 ( .IN(n6479), .QN(n6298) );
  INVX0 U5522 ( .IN(n6483), .QN(n6291) );
  INVX0 U5523 ( .IN(n6487), .QN(n6282) );
  INVX0 U5524 ( .IN(n6480), .QN(n6297) );
  INVX0 U5525 ( .IN(n6482), .QN(n6293) );
  INVX0 U5526 ( .IN(n6486), .QN(n6285) );
  INVX0 U5527 ( .IN(n6481), .QN(n6294) );
  INVX0 U5528 ( .IN(n6485), .QN(n6286) );
  INVX0 U5529 ( .IN(n6488), .QN(n6280) );
  INVX0 U5530 ( .IN(n6488), .QN(n6281) );
  INVX0 U5531 ( .IN(n6482), .QN(n6292) );
  INVX0 U5532 ( .IN(n6480), .QN(n6296) );
  INVX0 U5533 ( .IN(n6487), .QN(n6283) );
  INVX0 U5534 ( .IN(n6489), .QN(n6278) );
  INVX0 U5535 ( .IN(n6486), .QN(n6284) );
  INVX0 U5536 ( .IN(n6490), .QN(n6277) );
  INVX0 U5537 ( .IN(n6479), .QN(n6299) );
  INVX0 U5538 ( .IN(n6478), .QN(n6300) );
  INVX0 U5539 ( .IN(n6476), .QN(n6304) );
  INVX0 U5540 ( .IN(n6474), .QN(n6308) );
  INVX0 U5541 ( .IN(n6475), .QN(n6307) );
  INVX0 U5542 ( .IN(n6469), .QN(n6318) );
  INVX0 U5543 ( .IN(n6467), .QN(n6323) );
  INVX0 U5544 ( .IN(n6476), .QN(n6305) );
  INVX0 U5545 ( .IN(n6475), .QN(n6306) );
  INVX0 U5546 ( .IN(n6474), .QN(n6309) );
  INVX0 U5547 ( .IN(n6472), .QN(n6312) );
  INVX0 U5548 ( .IN(n6473), .QN(n6310) );
  INVX0 U5549 ( .IN(n6470), .QN(n6316) );
  INVX0 U5550 ( .IN(n6467), .QN(n6322) );
  INVX0 U5551 ( .IN(n6469), .QN(n6319) );
  INVX0 U5552 ( .IN(n6477), .QN(n6302) );
  INVX0 U5553 ( .IN(n6473), .QN(n6311) );
  INVX0 U5554 ( .IN(n6468), .QN(n6321) );
  INVX0 U5555 ( .IN(n6468), .QN(n6320) );
  INVX0 U5556 ( .IN(n6471), .QN(n6314) );
  INVX0 U5557 ( .IN(n6470), .QN(n6317) );
  INVX0 U5558 ( .IN(n6477), .QN(n6303) );
  INVX0 U5559 ( .IN(n6478), .QN(n6301) );
  INVX0 U5560 ( .IN(n6471), .QN(n6315) );
  INVX0 U5561 ( .IN(n6472), .QN(n6313) );
  INVX0 U5562 ( .IN(n6466), .QN(n6324) );
  INVX0 U5563 ( .IN(n6465), .QN(n6326) );
  INVX0 U5564 ( .IN(n6466), .QN(n6325) );
  INVX0 U5565 ( .IN(n6455), .QN(n6347) );
  INVX0 U5566 ( .IN(n6465), .QN(n6327) );
  INVX0 U5567 ( .IN(n6462), .QN(n6332) );
  INVX0 U5568 ( .IN(n6456), .QN(n6345) );
  INVX0 U5569 ( .IN(n6457), .QN(n6343) );
  INVX0 U5570 ( .IN(n6460), .QN(n6337) );
  INVX0 U5571 ( .IN(n6454), .QN(n6348) );
  INVX0 U5572 ( .IN(n6462), .QN(n6333) );
  INVX0 U5573 ( .IN(n6461), .QN(n6335) );
  INVX0 U5574 ( .IN(n6453), .QN(n6351) );
  INVX0 U5575 ( .IN(n6459), .QN(n6339) );
  INVX0 U5576 ( .IN(n6461), .QN(n6334) );
  INVX0 U5577 ( .IN(n6455), .QN(n6346) );
  INVX0 U5578 ( .IN(n6456), .QN(n6344) );
  INVX0 U5579 ( .IN(n6463), .QN(n6330) );
  INVX0 U5580 ( .IN(n6460), .QN(n6336) );
  INVX0 U5581 ( .IN(n6464), .QN(n6329) );
  INVX0 U5582 ( .IN(n6454), .QN(n6349) );
  INVX0 U5583 ( .IN(n6464), .QN(n6328) );
  INVX0 U5584 ( .IN(n6457), .QN(n6342) );
  INVX0 U5585 ( .IN(n6459), .QN(n6338) );
  INVX0 U5586 ( .IN(n6458), .QN(n6340) );
  INVX0 U5587 ( .IN(n6463), .QN(n6331) );
  INVX0 U5588 ( .IN(n6458), .QN(n6341) );
  INVX0 U5589 ( .IN(n6453), .QN(n6350) );
  INVX0 U5590 ( .IN(n6452), .QN(n6352) );
  INVX0 U5591 ( .IN(n6441), .QN(n6374) );
  INVX0 U5592 ( .IN(n6436), .QN(n6385) );
  INVX0 U5593 ( .IN(n6438), .QN(n6381) );
  INVX0 U5594 ( .IN(n6437), .QN(n6383) );
  INVX0 U5595 ( .IN(n6443), .QN(n6371) );
  INVX0 U5596 ( .IN(n6432), .QN(n6393) );
  INVX0 U5597 ( .IN(n6445), .QN(n6366) );
  INVX0 U5598 ( .IN(n6444), .QN(n6368) );
  INVX0 U5599 ( .IN(n6446), .QN(n6364) );
  INVX0 U5600 ( .IN(n6449), .QN(n6358) );
  INVX0 U5601 ( .IN(n6448), .QN(n6361) );
  INVX0 U5602 ( .IN(n6439), .QN(n6379) );
  INVX0 U5603 ( .IN(n6435), .QN(n6387) );
  INVX0 U5604 ( .IN(n6445), .QN(n6367) );
  INVX0 U5605 ( .IN(n6437), .QN(n6382) );
  INVX0 U5606 ( .IN(n6431), .QN(n6394) );
  INVX0 U5607 ( .IN(n6431), .QN(n6395) );
  INVX0 U5608 ( .IN(n6450), .QN(n6356) );
  INVX0 U5609 ( .IN(n6443), .QN(n6370) );
  INVX0 U5610 ( .IN(n6449), .QN(n6359) );
  INVX0 U5611 ( .IN(n6446), .QN(n6365) );
  INVX0 U5612 ( .IN(n6438), .QN(n6380) );
  INVX0 U5613 ( .IN(n6451), .QN(n6354) );
  INVX0 U5614 ( .IN(n6447), .QN(n6362) );
  INVX0 U5615 ( .IN(n6451), .QN(n6355) );
  INVX0 U5616 ( .IN(n6447), .QN(n6363) );
  INVX0 U5617 ( .IN(n6432), .QN(n6392) );
  INVX0 U5618 ( .IN(n6435), .QN(n6386) );
  INVX0 U5619 ( .IN(n6430), .QN(n6396) );
  INVX0 U5620 ( .IN(n6441), .QN(n6375) );
  INVX0 U5621 ( .IN(n6440), .QN(n6376) );
  INVX0 U5622 ( .IN(n6439), .QN(n6378) );
  INVX0 U5623 ( .IN(n6430), .QN(n6397) );
  INVX0 U5624 ( .IN(n6440), .QN(n6377) );
  INVX0 U5625 ( .IN(n6434), .QN(n6389) );
  INVX0 U5626 ( .IN(n6433), .QN(n6391) );
  INVX0 U5627 ( .IN(n6434), .QN(n6388) );
  INVX0 U5628 ( .IN(n6433), .QN(n6390) );
  INVX0 U5629 ( .IN(n6436), .QN(n6384) );
  INVX0 U5630 ( .IN(n6442), .QN(n6373) );
  INVX0 U5631 ( .IN(n6444), .QN(n6369) );
  INVX0 U5632 ( .IN(n6547), .QN(n6158) );
  INVX0 U5633 ( .IN(n6546), .QN(n6160) );
  INVX0 U5634 ( .IN(n6544), .QN(n6164) );
  INVX0 U5635 ( .IN(n6540), .QN(n6172) );
  INVX0 U5636 ( .IN(n6603), .QN(n6452) );
  INVX0 U5637 ( .IN(n6582), .QN(n6495) );
  INVX0 U5638 ( .IN(n6581), .QN(n6497) );
  INVX0 U5639 ( .IN(n6605), .QN(n6448) );
  INVX0 U5640 ( .IN(n6604), .QN(n6450) );
  INVX0 U5641 ( .IN(n6574), .QN(n6510) );
  INVX0 U5642 ( .IN(n6608), .QN(n6442) );
  INVX0 U5643 ( .IN(n6546), .QN(n6159) );
  INVX0 U5644 ( .IN(n6550), .QN(n6152) );
  INVX0 U5645 ( .IN(n6551), .QN(n6150) );
  INVX0 U5646 ( .IN(n6552), .QN(n6148) );
  INVX0 U5647 ( .IN(n6544), .QN(n6163) );
  INVX0 U5648 ( .IN(n6548), .QN(n6156) );
  INVX0 U5649 ( .IN(n6547), .QN(n6157) );
  INVX0 U5650 ( .IN(n6549), .QN(n6153) );
  INVX0 U5651 ( .IN(n6545), .QN(n6161) );
  INVX0 U5652 ( .IN(n6552), .QN(n6147) );
  INVX0 U5653 ( .IN(n6545), .QN(n6162) );
  INVX0 U5654 ( .IN(n6550), .QN(n6151) );
  INVX0 U5655 ( .IN(n6548), .QN(n6155) );
  INVX0 U5656 ( .IN(n6549), .QN(n6154) );
  INVX0 U5657 ( .IN(n6551), .QN(n6149) );
  INVX0 U5658 ( .IN(n6543), .QN(n6165) );
  INVX0 U5659 ( .IN(n6542), .QN(n6167) );
  INVX0 U5660 ( .IN(n6543), .QN(n6166) );
  INVX0 U5661 ( .IN(n6539), .QN(n6174) );
  INVX0 U5662 ( .IN(n6541), .QN(n6169) );
  INVX0 U5663 ( .IN(n6542), .QN(n6168) );
  INVX0 U5664 ( .IN(n6539), .QN(n6173) );
  INVX0 U5665 ( .IN(n6538), .QN(n6176) );
  INVX0 U5666 ( .IN(n6541), .QN(n6170) );
  INVX0 U5667 ( .IN(n6540), .QN(n6171) );
  INVX0 U5668 ( .IN(n6538), .QN(n6175) );
  INVX0 U5669 ( .IN(n6537), .QN(n6177) );
  INVX0 U5670 ( .IN(n6537), .QN(n6178) );
  INVX0 U5671 ( .IN(n6536), .QN(n6180) );
  INVX0 U5672 ( .IN(n6536), .QN(n6179) );
  INVX0 U5673 ( .IN(n6533), .QN(n6186) );
  INVX0 U5674 ( .IN(n6533), .QN(n6185) );
  INVX0 U5675 ( .IN(n6534), .QN(n6183) );
  INVX0 U5676 ( .IN(n6532), .QN(n6188) );
  INVX0 U5677 ( .IN(n6531), .QN(n6189) );
  INVX0 U5678 ( .IN(n6532), .QN(n6187) );
  INVX0 U5679 ( .IN(n6534), .QN(n6184) );
  INVX0 U5680 ( .IN(n6529), .QN(n6194) );
  INVX0 U5681 ( .IN(n6530), .QN(n6192) );
  INVX0 U5682 ( .IN(n6535), .QN(n6181) );
  INVX0 U5683 ( .IN(n6529), .QN(n6193) );
  INVX0 U5684 ( .IN(n6531), .QN(n6190) );
  INVX0 U5685 ( .IN(n6530), .QN(n6191) );
  INVX0 U5686 ( .IN(n6535), .QN(n6182) );
  INVX0 U5687 ( .IN(n6528), .QN(n6195) );
  INVX0 U5688 ( .IN(n6527), .QN(n6198) );
  INVX0 U5689 ( .IN(n6527), .QN(n6197) );
  INVX0 U5690 ( .IN(n6528), .QN(n6196) );
  INVX0 U5691 ( .IN(n6525), .QN(n6201) );
  INVX0 U5692 ( .IN(n6525), .QN(n6202) );
  INVX0 U5693 ( .IN(n6526), .QN(n6200) );
  INVX0 U5694 ( .IN(n6526), .QN(n6199) );
  INVX0 U5695 ( .IN(n6524), .QN(n6203) );
  INVX0 U5696 ( .IN(n6524), .QN(n6204) );
  INVX0 U5697 ( .IN(n6522), .QN(n6208) );
  INVX0 U5698 ( .IN(n6523), .QN(n6205) );
  INVX0 U5699 ( .IN(n6521), .QN(n6209) );
  INVX0 U5700 ( .IN(n6521), .QN(n6210) );
  INVX0 U5701 ( .IN(n6523), .QN(n6206) );
  INVX0 U5702 ( .IN(n6522), .QN(n6207) );
  INVX0 U5703 ( .IN(n6424), .QN(n6409) );
  INVX0 U5704 ( .IN(n6426), .QN(n6404) );
  INVX0 U5705 ( .IN(n6422), .QN(n6413) );
  INVX0 U5706 ( .IN(n6422), .QN(n6412) );
  INVX0 U5707 ( .IN(n6428), .QN(n6400) );
  INVX0 U5708 ( .IN(n6425), .QN(n6407) );
  INVX0 U5709 ( .IN(n6426), .QN(n6405) );
  INVX0 U5710 ( .IN(n6427), .QN(n6402) );
  INVX0 U5711 ( .IN(n6427), .QN(n6403) );
  INVX0 U5712 ( .IN(n6429), .QN(n6399) );
  INVX0 U5713 ( .IN(n6428), .QN(n6401) );
  INVX0 U5714 ( .IN(n6423), .QN(n6411) );
  INVX0 U5715 ( .IN(n6423), .QN(n6410) );
  INVX0 U5716 ( .IN(n6429), .QN(n6398) );
  INVX0 U5717 ( .IN(n6424), .QN(n6408) );
  INVX0 U5718 ( .IN(n6425), .QN(n6406) );
  INVX0 U5719 ( .IN(n6581), .QN(n6496) );
  INVX0 U5720 ( .IN(n6577), .QN(n6504) );
  INVX0 U5721 ( .IN(n6569), .QN(n6520) );
  INVX0 U5722 ( .IN(n6569), .QN(n6519) );
  INVX0 U5723 ( .IN(n6573), .QN(n6513) );
  INVX0 U5724 ( .IN(n6607), .QN(n6444) );
  INVX0 U5725 ( .IN(n6570), .QN(n6517) );
  INVX0 U5726 ( .IN(n6607), .QN(n6445) );
  INVX0 U5727 ( .IN(n6611), .QN(n6437) );
  INVX0 U5728 ( .IN(n6614), .QN(n6431) );
  INVX0 U5729 ( .IN(n6608), .QN(n6443) );
  INVX0 U5730 ( .IN(n6605), .QN(n6449) );
  INVX0 U5731 ( .IN(n6606), .QN(n6446) );
  INVX0 U5732 ( .IN(n6610), .QN(n6438) );
  INVX0 U5733 ( .IN(n6665), .QN(n6511) );
  INVX0 U5734 ( .IN(n6604), .QN(n6451) );
  INVX0 U5735 ( .IN(n6606), .QN(n6447) );
  INVX0 U5736 ( .IN(n6572), .QN(n6515) );
  INVX0 U5737 ( .IN(n6613), .QN(n6432) );
  INVX0 U5738 ( .IN(n6612), .QN(n6435) );
  INVX0 U5739 ( .IN(n6570), .QN(n6518) );
  INVX0 U5740 ( .IN(n6572), .QN(n6516) );
  INVX0 U5741 ( .IN(n6609), .QN(n6441) );
  INVX0 U5742 ( .IN(n6610), .QN(n6439) );
  INVX0 U5743 ( .IN(n6573), .QN(n6514) );
  INVX0 U5744 ( .IN(n6614), .QN(n6430) );
  INVX0 U5745 ( .IN(n6609), .QN(n6440) );
  INVX0 U5746 ( .IN(n6597), .QN(n6465) );
  INVX0 U5747 ( .IN(n6575), .QN(n6508) );
  INVX0 U5748 ( .IN(n6612), .QN(n6434) );
  INVX0 U5749 ( .IN(n6613), .QN(n6433) );
  INVX0 U5750 ( .IN(n6576), .QN(n6507) );
  INVX0 U5751 ( .IN(n6668), .QN(n6512) );
  INVX0 U5752 ( .IN(n6577), .QN(n6505) );
  INVX0 U5753 ( .IN(n6596), .QN(n6466) );
  INVX0 U5754 ( .IN(n6579), .QN(n6501) );
  INVX0 U5755 ( .IN(n6578), .QN(n6502) );
  INVX0 U5756 ( .IN(n6611), .QN(n6436) );
  INVX0 U5757 ( .IN(n6578), .QN(n6503) );
  INVX0 U5758 ( .IN(n6576), .QN(n6506) );
  INVX0 U5759 ( .IN(n6579), .QN(n6500) );
  INVX0 U5760 ( .IN(n6575), .QN(n6509) );
  INVX0 U5761 ( .IN(n6580), .QN(n6499) );
  INVX0 U5762 ( .IN(n6591), .QN(n6476) );
  INVX0 U5763 ( .IN(n6592), .QN(n6475) );
  INVX0 U5764 ( .IN(n6598), .QN(n6462) );
  INVX0 U5765 ( .IN(n6587), .QN(n6484) );
  INVX0 U5766 ( .IN(n6592), .QN(n6474) );
  INVX0 U5767 ( .IN(n6599), .QN(n6461) );
  INVX0 U5768 ( .IN(n6596), .QN(n6467) );
  INVX0 U5769 ( .IN(n6602), .QN(n6455) );
  INVX0 U5770 ( .IN(n6590), .QN(n6479) );
  INVX0 U5771 ( .IN(n6588), .QN(n6483) );
  INVX0 U5772 ( .IN(n6601), .QN(n6456) );
  INVX0 U5773 ( .IN(n6589), .QN(n6481) );
  INVX0 U5774 ( .IN(n6599), .QN(n6460) );
  INVX0 U5775 ( .IN(n6595), .QN(n6469) );
  INVX0 U5776 ( .IN(n6593), .QN(n6473) );
  INVX0 U5777 ( .IN(n6602), .QN(n6454) );
  INVX0 U5778 ( .IN(n6595), .QN(n6468) );
  INVX0 U5779 ( .IN(n6587), .QN(n6485) );
  INVX0 U5780 ( .IN(n6597), .QN(n6464) );
  INVX0 U5781 ( .IN(n6582), .QN(n6494) );
  INVX0 U5782 ( .IN(n6583), .QN(n6492) );
  INVX0 U5783 ( .IN(n6594), .QN(n6470) );
  INVX0 U5784 ( .IN(n6585), .QN(n6488) );
  INVX0 U5785 ( .IN(n6601), .QN(n6457) );
  INVX0 U5786 ( .IN(n6591), .QN(n6477) );
  INVX0 U5787 ( .IN(n6588), .QN(n6482) );
  INVX0 U5788 ( .IN(n6589), .QN(n6480) );
  INVX0 U5789 ( .IN(n6586), .QN(n6487) );
  INVX0 U5790 ( .IN(n6583), .QN(n6493) );
  INVX0 U5791 ( .IN(n6585), .QN(n6489) );
  INVX0 U5792 ( .IN(n6600), .QN(n6459) );
  INVX0 U5793 ( .IN(n6586), .QN(n6486) );
  INVX0 U5794 ( .IN(n6598), .QN(n6463) );
  INVX0 U5795 ( .IN(n6584), .QN(n6490) );
  INVX0 U5796 ( .IN(n6590), .QN(n6478) );
  INVX0 U5797 ( .IN(n6600), .QN(n6458) );
  INVX0 U5798 ( .IN(n6584), .QN(n6491) );
  INVX0 U5799 ( .IN(n6594), .QN(n6471) );
  INVX0 U5800 ( .IN(n6603), .QN(n6453) );
  INVX0 U5801 ( .IN(n6593), .QN(n6472) );
  INVX0 U5802 ( .IN(n6639), .QN(n6580) );
  INVX0 U5803 ( .IN(n6555), .QN(n6547) );
  INVX0 U5804 ( .IN(n6556), .QN(n6546) );
  INVX0 U5805 ( .IN(n6557), .QN(n6544) );
  INVX0 U5806 ( .IN(n6627), .QN(n6603) );
  INVX0 U5807 ( .IN(n6638), .QN(n6582) );
  INVX0 U5808 ( .IN(n6638), .QN(n6581) );
  INVX0 U5809 ( .IN(n6626), .QN(n6605) );
  INVX0 U5810 ( .IN(n6627), .QN(n6604) );
  INVX0 U5811 ( .IN(n6642), .QN(n6574) );
  INVX0 U5812 ( .IN(n6625), .QN(n6608) );
  INVX0 U5813 ( .IN(n6559), .QN(n6540) );
  INVX0 U5814 ( .IN(n6421), .QN(n6414) );
  INVX0 U5815 ( .IN(n6420), .QN(n6417) );
  INVX0 U5816 ( .IN(n6421), .QN(n6415) );
  INVX0 U5817 ( .IN(n6420), .QN(n6416) );
  INVX0 U5818 ( .IN(n6640), .QN(n6577) );
  INVX0 U5819 ( .IN(n6644), .QN(n6569) );
  INVX0 U5820 ( .IN(n6554), .QN(n6550) );
  INVX0 U5821 ( .IN(n6553), .QN(n6551) );
  INVX0 U5822 ( .IN(n6553), .QN(n6552) );
  INVX0 U5823 ( .IN(n6560), .QN(n6537) );
  INVX0 U5824 ( .IN(n6625), .QN(n6607) );
  INVX0 U5825 ( .IN(n6558), .QN(n6542) );
  INVX0 U5826 ( .IN(n6557), .QN(n6543) );
  INVX0 U5827 ( .IN(n6626), .QN(n6606) );
  INVX0 U5828 ( .IN(n6644), .QN(n6570) );
  INVX0 U5829 ( .IN(n6643), .QN(n6572) );
  INVX0 U5830 ( .IN(n6624), .QN(n6610) );
  INVX0 U5831 ( .IN(n6673), .QN(n6573) );
  INVX0 U5832 ( .IN(n6622), .QN(n6614) );
  INVX0 U5833 ( .IN(n6643), .QN(n6571) );
  INVX0 U5834 ( .IN(n6624), .QN(n6609) );
  INVX0 U5835 ( .IN(n6630), .QN(n6597) );
  INVX0 U5836 ( .IN(n6555), .QN(n6548) );
  INVX0 U5837 ( .IN(n6623), .QN(n6612) );
  INVX0 U5838 ( .IN(n6622), .QN(n6613) );
  INVX0 U5839 ( .IN(n6631), .QN(n6596) );
  INVX0 U5840 ( .IN(n6623), .QN(n6611) );
  INVX0 U5841 ( .IN(n6640), .QN(n6578) );
  INVX0 U5842 ( .IN(n6641), .QN(n6576) );
  INVX0 U5843 ( .IN(n6639), .QN(n6579) );
  INVX0 U5844 ( .IN(n6641), .QN(n6575) );
  INVX0 U5845 ( .IN(n6554), .QN(n6549) );
  INVX0 U5846 ( .IN(n6562), .QN(n6533) );
  INVX0 U5847 ( .IN(n6559), .QN(n6539) );
  INVX0 U5848 ( .IN(n6556), .QN(n6545) );
  INVX0 U5849 ( .IN(n6618), .QN(n6422) );
  INVX0 U5850 ( .IN(n6558), .QN(n6541) );
  INVX0 U5851 ( .IN(n6563), .QN(n6532) );
  INVX0 U5852 ( .IN(n6616), .QN(n6426) );
  INVX0 U5853 ( .IN(n6562), .QN(n6534) );
  INVX0 U5854 ( .IN(n6633), .QN(n6592) );
  INVX0 U5855 ( .IN(n6616), .QN(n6427) );
  INVX0 U5856 ( .IN(n6567), .QN(n6524) );
  INVX0 U5857 ( .IN(n6568), .QN(n6521) );
  INVX0 U5858 ( .IN(n6565), .QN(n6527) );
  INVX0 U5859 ( .IN(n6615), .QN(n6428) );
  INVX0 U5860 ( .IN(n6567), .QN(n6523) );
  INVX0 U5861 ( .IN(n6565), .QN(n6528) );
  INVX0 U5862 ( .IN(n6629), .QN(n6599) );
  INVX0 U5863 ( .IN(n6566), .QN(n6525) );
  INVX0 U5864 ( .IN(n6561), .QN(n6536) );
  INVX0 U5865 ( .IN(n6566), .QN(n6526) );
  INVX0 U5866 ( .IN(n6628), .QN(n6602) );
  INVX0 U5867 ( .IN(n6631), .QN(n6595) );
  INVX0 U5868 ( .IN(n6635), .QN(n6587) );
  INVX0 U5869 ( .IN(n6564), .QN(n6529) );
  INVX0 U5870 ( .IN(n6628), .QN(n6601) );
  INVX0 U5871 ( .IN(n6633), .QN(n6591) );
  INVX0 U5872 ( .IN(n6560), .QN(n6538) );
  INVX0 U5873 ( .IN(n6618), .QN(n6423) );
  INVX0 U5874 ( .IN(n6635), .QN(n6588) );
  INVX0 U5875 ( .IN(n6634), .QN(n6589) );
  INVX0 U5876 ( .IN(n6615), .QN(n6429) );
  INVX0 U5877 ( .IN(n6617), .QN(n6424) );
  INVX0 U5878 ( .IN(n6637), .QN(n6583) );
  INVX0 U5879 ( .IN(n6636), .QN(n6585) );
  INVX0 U5880 ( .IN(n6636), .QN(n6586) );
  INVX0 U5881 ( .IN(n6630), .QN(n6598) );
  INVX0 U5882 ( .IN(n6634), .QN(n6590) );
  INVX0 U5883 ( .IN(n6629), .QN(n6600) );
  INVX0 U5884 ( .IN(n6637), .QN(n6584) );
  INVX0 U5885 ( .IN(n6563), .QN(n6531) );
  INVX0 U5886 ( .IN(n6617), .QN(n6425) );
  INVX0 U5887 ( .IN(n6632), .QN(n6594) );
  INVX0 U5888 ( .IN(n6568), .QN(n6522) );
  INVX0 U5889 ( .IN(n6564), .QN(n6530) );
  INVX0 U5890 ( .IN(n6561), .QN(n6535) );
  INVX0 U5891 ( .IN(n6632), .QN(n6593) );
  INVX0 U5892 ( .IN(n6651), .QN(n6555) );
  INVX0 U5893 ( .IN(n6651), .QN(n6556) );
  INVX0 U5894 ( .IN(n6650), .QN(n6557) );
  INVX0 U5895 ( .IN(n6666), .QN(n6627) );
  INVX0 U5896 ( .IN(n6660), .QN(n6638) );
  INVX0 U5897 ( .IN(n6666), .QN(n6626) );
  INVX0 U5898 ( .IN(n6658), .QN(n6642) );
  INVX0 U5899 ( .IN(n6667), .QN(n6625) );
  INVX0 U5900 ( .IN(n6649), .QN(n6559) );
  NBUFFX2 U5901 ( .IN(n6057), .Q(n6029) );
  NBUFFX2 U5902 ( .IN(n6056), .Q(n6031) );
  NBUFFX2 U5903 ( .IN(n6055), .Q(n6033) );
  NBUFFX2 U5904 ( .IN(n6056), .Q(n6032) );
  NBUFFX2 U5905 ( .IN(n6055), .Q(n6034) );
  NBUFFX2 U5906 ( .IN(n6057), .Q(n6030) );
  NBUFFX2 U5907 ( .IN(n6054), .Q(n6035) );
  NBUFFX2 U5908 ( .IN(n6054), .Q(n6036) );
  NBUFFX2 U5909 ( .IN(n6050), .Q(n6044) );
  NBUFFX2 U5910 ( .IN(n6051), .Q(n6041) );
  NBUFFX2 U5911 ( .IN(n6052), .Q(n6040) );
  NBUFFX2 U5912 ( .IN(n6052), .Q(n6039) );
  NBUFFX2 U5913 ( .IN(n6049), .Q(n6045) );
  NBUFFX2 U5914 ( .IN(n6051), .Q(n6042) );
  NBUFFX2 U5915 ( .IN(n6053), .Q(n6037) );
  NBUFFX2 U5916 ( .IN(n6050), .Q(n6043) );
  NBUFFX2 U5917 ( .IN(n6053), .Q(n6038) );
  NBUFFX2 U5918 ( .IN(n6049), .Q(n6046) );
  INVX0 U5919 ( .IN(n6633), .QN(n6418) );
  INVX0 U5920 ( .IN(n6659), .QN(n6640) );
  INVX0 U5921 ( .IN(n6657), .QN(n6644) );
  INVX0 U5922 ( .IN(n6652), .QN(n6553) );
  INVX0 U5923 ( .IN(n6649), .QN(n6560) );
  INVX0 U5924 ( .IN(n6650), .QN(n6558) );
  INVX0 U5925 ( .IN(n6657), .QN(n6643) );
  INVX0 U5926 ( .IN(n6667), .QN(n6624) );
  INVX0 U5927 ( .IN(n6664), .QN(n6630) );
  INVX0 U5928 ( .IN(n6668), .QN(n6622) );
  INVX0 U5929 ( .IN(n6664), .QN(n6631) );
  INVX0 U5930 ( .IN(n6668), .QN(n6623) );
  INVX0 U5931 ( .IN(n6659), .QN(n6641) );
  INVX0 U5932 ( .IN(n6652), .QN(n6554) );
  INVX0 U5933 ( .IN(n6619), .QN(n6420) );
  INVX0 U5934 ( .IN(n6648), .QN(n6562) );
  INVX0 U5935 ( .IN(n6621), .QN(n6616) );
  INVX0 U5936 ( .IN(n6645), .QN(n6567) );
  INVX0 U5937 ( .IN(n6646), .QN(n6565) );
  INVX0 U5938 ( .IN(n6646), .QN(n6566) );
  INVX0 U5939 ( .IN(n6619), .QN(n6421) );
  INVX0 U5940 ( .IN(n6665), .QN(n6628) );
  INVX0 U5941 ( .IN(n6663), .QN(n6633) );
  INVX0 U5942 ( .IN(n6620), .QN(n6618) );
  INVX0 U5943 ( .IN(n6662), .QN(n6635) );
  INVX0 U5944 ( .IN(n6621), .QN(n6615) );
  INVX0 U5945 ( .IN(n6661), .QN(n6636) );
  INVX0 U5946 ( .IN(n6662), .QN(n6634) );
  INVX0 U5947 ( .IN(n6665), .QN(n6629) );
  INVX0 U5948 ( .IN(n6661), .QN(n6637) );
  INVX0 U5949 ( .IN(n6647), .QN(n6563) );
  INVX0 U5950 ( .IN(n6620), .QN(n6617) );
  INVX0 U5951 ( .IN(n6645), .QN(n6568) );
  INVX0 U5952 ( .IN(n6647), .QN(n6564) );
  INVX0 U5953 ( .IN(n6648), .QN(n6561) );
  INVX0 U5954 ( .IN(n6663), .QN(n6632) );
  INVX0 U5955 ( .IN(n6637), .QN(n6419) );
  NBUFFX2 U5956 ( .IN(n6048), .Q(n6047) );
  INVX0 U5957 ( .IN(n2748), .QN(n1305) );
  INVX0 U5958 ( .IN(n2763), .QN(n1301) );
  INVX0 U5959 ( .IN(n3498), .QN(n1279) );
  INVX0 U5960 ( .IN(n6674), .QN(n6660) );
  ISOLANDX1 U5961 ( .D(n3593), .ISO(n3589), .Q(n3595) );
  ISOLANDX1 U5962 ( .D(n3574), .ISO(n3570), .Q(n3576) );
  ISOLANDX1 U5963 ( .D(n3517), .ISO(n3513), .Q(n3519) );
  ISOLANDX1 U5964 ( .D(n3628), .ISO(n3624), .Q(n3630) );
  ISOLANDX1 U5965 ( .D(n3555), .ISO(n3551), .Q(n3557) );
  ISOLANDX1 U5966 ( .D(n3646), .ISO(n3642), .Q(n3648) );
  ISOLANDX1 U5967 ( .D(n3536), .ISO(n3532), .Q(n3538) );
  ISOLANDX1 U5968 ( .D(n3611), .ISO(n3607), .Q(n3613) );
  INVX0 U5969 ( .IN(n6653), .QN(n6651) );
  INVX0 U5970 ( .IN(n6654), .QN(n6650) );
  INVX0 U5971 ( .IN(n6671), .QN(n6666) );
  INVX0 U5972 ( .IN(n6654), .QN(n6649) );
  INVX0 U5973 ( .IN(n6675), .QN(n6658) );
  INVX0 U5974 ( .IN(n6670), .QN(n6667) );
  NAND2X0 U5975 ( .IN1(n1461), .IN2(n6080), .QN(n3305) );
  NBUFFX2 U5976 ( .IN(n6058), .Q(n6056) );
  NBUFFX2 U5977 ( .IN(n6059), .Q(n6055) );
  NBUFFX2 U5978 ( .IN(n6058), .Q(n6057) );
  NBUFFX2 U5979 ( .IN(n6059), .Q(n6054) );
  NBUFFX2 U5980 ( .IN(n6060), .Q(n6052) );
  NBUFFX2 U5981 ( .IN(n6062), .Q(n6049) );
  NBUFFX2 U5982 ( .IN(n6061), .Q(n6051) );
  NBUFFX2 U5983 ( .IN(n6061), .Q(n6050) );
  NBUFFX2 U5984 ( .IN(n6060), .Q(n6053) );
  INVX0 U5985 ( .IN(n2688), .QN(n1554) );
  INVX0 U5986 ( .IN(n2667), .QN(n1700) );
  NAND2X0 U5987 ( .IN1(n1306), .IN2(n6178), .QN(n2748) );
  NAND2X0 U5988 ( .IN1(n1302), .IN2(n6179), .QN(n2763) );
  NAND2X0 U5989 ( .IN1(n6198), .IN2(n3503), .QN(n3498) );
  INVX0 U5990 ( .IN(n4545), .QN(n1449) );
  NOR2X0 U5991 ( .IN1(n2966), .IN2(n6067), .QN(n2957) );
  NOR2X0 U5992 ( .IN1(n2906), .IN2(n6067), .QN(n2887) );
  NOR2X0 U5993 ( .IN1(n2930), .IN2(n6067), .QN(n2911) );
  NOR2X0 U5994 ( .IN1(n2953), .IN2(n6067), .QN(n2934) );
  NOR2X0 U5995 ( .IN1(n1337), .IN2(n6066), .QN(n2793) );
  NOR2X0 U5996 ( .IN1(n1313), .IN2(n6066), .QN(n2863) );
  NOR2X0 U5997 ( .IN1(n1329), .IN2(n6066), .QN(n2817) );
  NOR2X0 U5998 ( .IN1(n1321), .IN2(n6066), .QN(n2840) );
  INVX0 U5999 ( .IN(n6674), .QN(n6659) );
  INVX0 U6000 ( .IN(n6675), .QN(n6657) );
  INVX0 U6001 ( .IN(n6672), .QN(n6664) );
  INVX0 U6002 ( .IN(n6670), .QN(n6668) );
  INVX0 U6003 ( .IN(n6653), .QN(n6652) );
  INVX0 U6004 ( .IN(n6656), .QN(n6646) );
  INVX0 U6005 ( .IN(n6673), .QN(n6619) );
  INVX0 U6006 ( .IN(n6669), .QN(n6621) );
  INVX0 U6007 ( .IN(n6673), .QN(n6662) );
  INVX0 U6008 ( .IN(n6671), .QN(n6665) );
  INVX0 U6009 ( .IN(n6673), .QN(n6661) );
  INVX0 U6010 ( .IN(n6669), .QN(n6620) );
  INVX0 U6011 ( .IN(n6656), .QN(n6645) );
  INVX0 U6012 ( .IN(n6655), .QN(n6647) );
  INVX0 U6013 ( .IN(n6655), .QN(n6648) );
  INVX0 U6014 ( .IN(n6672), .QN(n6663) );
  NAND2X0 U6015 ( .IN1(n1298), .IN2(n6163), .QN(n2587) );
  NOR2X0 U6016 ( .IN1(n1469), .IN2(n1470), .QN(n3008) );
  NBUFFX2 U6017 ( .IN(n6062), .Q(n6048) );
  INVX0 U6018 ( .IN(n3451), .QN(n1399) );
  INVX0 U6019 ( .IN(n2559), .QN(n1308) );
  INVX0 U6020 ( .IN(n2569), .QN(n1304) );
  INVX0 U6021 ( .IN(n2709), .QN(n1422) );
  INVX0 U6022 ( .IN(n3006), .QN(n1472) );
  INVX0 U6023 ( .IN(n3631), .QN(n1397) );
  INVX0 U6024 ( .IN(n3558), .QN(n1393) );
  INVX0 U6025 ( .IN(n3596), .QN(n1395) );
  INVX0 U6026 ( .IN(n3539), .QN(n1392) );
  INVX0 U6027 ( .IN(n3520), .QN(n1391) );
  INVX0 U6028 ( .IN(n3614), .QN(n1396) );
  INVX0 U6029 ( .IN(n3169), .QN(n1310) );
  INVX0 U6030 ( .IN(n3210), .QN(n1366) );
  INVX0 U6031 ( .IN(n3109), .QN(n1334) );
  INVX0 U6032 ( .IN(n3230), .QN(n1357) );
  INVX0 U6033 ( .IN(n3129), .QN(n1326) );
  INVX0 U6034 ( .IN(n3248), .QN(n1348) );
  INVX0 U6035 ( .IN(n3190), .QN(n1375) );
  INVX0 U6036 ( .IN(n3150), .QN(n1318) );
  INVX0 U6037 ( .IN(n3649), .QN(n1398) );
  INVX0 U6038 ( .IN(n3577), .QN(n1394) );
  INVX0 U6039 ( .IN(n2416), .QN(n1490) );
  INVX0 U6040 ( .IN(n5087), .QN(n1928) );
  INVX0 U6041 ( .IN(n3503), .QN(n1280) );
  INVX0 U6042 ( .IN(n3399), .QN(n1283) );
  INVX0 U6043 ( .IN(n3484), .QN(n1281) );
  INVX0 U6044 ( .IN(n3474), .QN(n1282) );
  INVX0 U6045 ( .IN(n4159), .QN(n1496) );
  AO21X1 U6046 ( .IN1(n3304), .IN2(n3352), .IN3(n3305), .Q(n3333) );
  NOR2X0 U6047 ( .IN1(n6083), .IN2(n1454), .QN(n2518) );
  NOR2X0 U6048 ( .IN1(n6082), .IN2(n1452), .QN(n2535) );
  NOR2X0 U6049 ( .IN1(n6082), .IN2(n1455), .QN(n2523) );
  NOR2X0 U6050 ( .IN1(n6082), .IN2(n1456), .QN(n2522) );
  NOR2X0 U6051 ( .IN1(n6082), .IN2(n1457), .QN(n2521) );
  NOR2X0 U6052 ( .IN1(n6080), .IN2(n1309), .QN(n2534) );
  NOR2X0 U6053 ( .IN1(n3627), .IN2(n6069), .QN(n3628) );
  NOR2X0 U6054 ( .IN1(n3554), .IN2(n6068), .QN(n3555) );
  NOR2X0 U6055 ( .IN1(n3592), .IN2(n6069), .QN(n3593) );
  NOR2X0 U6056 ( .IN1(n3516), .IN2(n6068), .QN(n3517) );
  NOR2X0 U6057 ( .IN1(n3535), .IN2(n6068), .QN(n3536) );
  NOR2X0 U6058 ( .IN1(n3610), .IN2(n6069), .QN(n3611) );
  NOR2X0 U6059 ( .IN1(n6081), .IN2(n1277), .QN(n2532) );
  NOR2X0 U6060 ( .IN1(n6081), .IN2(n1453), .QN(n2540) );
  INVX0 U6061 ( .IN(n6677), .QN(n6653) );
  INVX0 U6062 ( .IN(n6677), .QN(n6654) );
  INVX0 U6063 ( .IN(n6681), .QN(n6671) );
  INVX0 U6064 ( .IN(n6679), .QN(n6675) );
  INVX0 U6065 ( .IN(n6681), .QN(n6670) );
  NOR2X0 U6066 ( .IN1(n3645), .IN2(n6069), .QN(n3646) );
  NOR2X0 U6067 ( .IN1(n3573), .IN2(n6069), .QN(n3574) );
  NOR2X0 U6068 ( .IN1(n3757), .IN2(n1417), .QN(n2477) );
  NOR2X0 U6069 ( .IN1(n1277), .IN2(n2398), .QN(n2396) );
  NBUFFX2 U6070 ( .IN(n3765), .Q(n6059) );
  NBUFFX2 U6071 ( .IN(n3765), .Q(n6058) );
  NBUFFX2 U6072 ( .IN(n3765), .Q(n6062) );
  NBUFFX2 U6073 ( .IN(n3765), .Q(n6061) );
  NBUFFX2 U6074 ( .IN(n3765), .Q(n6060) );
  INVX0 U6075 ( .IN(n4842), .QN(n1424) );
  NAND2X0 U6076 ( .IN1(n6190), .IN2(n2076), .QN(n4545) );
  NOR2X0 U6077 ( .IN1(n2560), .IN2(n6078), .QN(n2559) );
  NOR2X0 U6078 ( .IN1(n2570), .IN2(n6077), .QN(n2569) );
  NAND2X0 U6079 ( .IN1(n6185), .IN2(n3627), .QN(n3631) );
  NAND2X0 U6080 ( .IN1(n6194), .IN2(n3554), .QN(n3558) );
  NAND2X0 U6081 ( .IN1(n1351), .IN2(n1599), .QN(n2966) );
  NAND2X0 U6082 ( .IN1(n6197), .IN2(n3592), .QN(n3596) );
  NAND2X0 U6083 ( .IN1(n6204), .IN2(n3516), .QN(n3520) );
  NAND2X0 U6084 ( .IN1(n6203), .IN2(n3535), .QN(n3539) );
  NAND2X0 U6085 ( .IN1(n6186), .IN2(n3610), .QN(n3614) );
  NAND2X0 U6086 ( .IN1(n3712), .IN2(n6153), .QN(n3451) );
  NAND2X0 U6087 ( .IN1(n2441), .IN2(n2442), .QN(g26875) );
  NAND2X0 U6088 ( .IN1(n3505), .IN2(n3525), .QN(n3006) );
  NAND2X0 U6089 ( .IN1(n1369), .IN2(n1602), .QN(n2930) );
  NAND2X0 U6090 ( .IN1(n1360), .IN2(n1601), .QN(n2953) );
  NAND2X0 U6091 ( .IN1(n1378), .IN2(n1600), .QN(n2906) );
  NAND2X0 U6092 ( .IN1(n1516), .IN2(n6162), .QN(n2709) );
  NOR2X0 U6093 ( .IN1(n3258), .IN2(n6067), .QN(n3658) );
  NOR2X0 U6094 ( .IN1(n3266), .IN2(n6067), .QN(n3667) );
  NAND2X0 U6095 ( .IN1(n6189), .IN2(n3645), .QN(n3649) );
  NAND2X0 U6096 ( .IN1(n6211), .IN2(n3573), .QN(n3577) );
  INVX0 U6097 ( .IN(n2615), .QN(n1288) );
  NAND2X0 U6098 ( .IN1(n1952), .IN2(n1855), .QN(n4145) );
  NAND2X0 U6099 ( .IN1(n1759), .IN2(n1745), .QN(n4097) );
  ISOLANDX1 U6100 ( .D(n3635), .ISO(n6145), .Q(n4888) );
  AND3X1 U6101 ( .IN1(n3315), .IN2(n3312), .IN3(n3314), .Q(n3304) );
  NOR2X0 U6102 ( .IN1(n3550), .IN2(n3554), .QN(n3553) );
  NOR2X0 U6103 ( .IN1(n1466), .IN2(n3627), .QN(n3626) );
  NOR2X0 U6104 ( .IN1(n6081), .IN2(n1611), .QN(n3072) );
  NOR2X0 U6105 ( .IN1(n6082), .IN2(n1565), .QN(n3030) );
  INVX0 U6106 ( .IN(n6680), .QN(n6672) );
  INVX0 U6107 ( .IN(n6680), .QN(n6673) );
  INVX0 U6108 ( .IN(n6672), .QN(n6669) );
  INVX0 U6109 ( .IN(n6676), .QN(n6656) );
  INVX0 U6110 ( .IN(n6676), .QN(n6655) );
  NOR2X0 U6111 ( .IN1(n2596), .IN2(n6079), .QN(n2595) );
  NAND3X0 U6112 ( .IN1(n2531), .IN2(n1461), .IN3(n2527), .QN(n3318) );
  NOR2X0 U6113 ( .IN1(n1560), .IN2(n6068), .QN(n3059) );
  NOR2X0 U6114 ( .IN1(n1562), .IN2(n6068), .QN(n3051) );
  NOR2X0 U6115 ( .IN1(n1590), .IN2(n6067), .QN(n3093) );
  NOR2X0 U6116 ( .IN1(n1705), .IN2(n6069), .QN(n3022) );
  NOR2X0 U6117 ( .IN1(n1564), .IN2(n6069), .QN(n3042) );
  NOR2X0 U6118 ( .IN1(n1650), .IN2(n6068), .QN(n3083) );
  NOR2X0 U6119 ( .IN1(n2615), .IN2(n1599), .QN(n3241) );
  INVX0 U6120 ( .IN(n3627), .QN(n1855) );
  INVX0 U6121 ( .IN(n3554), .QN(n1745) );
  NOR2X0 U6122 ( .IN1(n2612), .IN2(n6078), .QN(n2610) );
  NOR2X0 U6123 ( .IN1(n2626), .IN2(n6078), .QN(n2624) );
  NOR2X0 U6124 ( .IN1(n2622), .IN2(n6079), .QN(n2620) );
  NOR4X0 U6125 ( .IN1(n1474), .IN2(n1477), .IN3(n1479), .IN4(n1481), .QN(n2729) );
  INVX0 U6126 ( .IN(n6025), .QN(n1461) );
  NAND2X0 U6127 ( .IN1(n3524), .IN2(n3005), .QN(n3624) );
  INVX0 U6128 ( .IN(n2870), .QN(n1313) );
  INVX0 U6129 ( .IN(n2824), .QN(n1329) );
  INVX0 U6130 ( .IN(n2847), .QN(n1321) );
  INVX0 U6131 ( .IN(n2800), .QN(n1337) );
  NAND2X0 U6132 ( .IN1(n3524), .IN2(n1468), .QN(n3589) );
  NAND2X0 U6133 ( .IN1(n3524), .IN2(n1467), .QN(n3607) );
  NAND2X0 U6134 ( .IN1(n3524), .IN2(n1471), .QN(n3532) );
  NAND2X0 U6135 ( .IN1(n3524), .IN2(n1472), .QN(n3513) );
  NAND2X0 U6136 ( .IN1(n3524), .IN2(n1469), .QN(n3570) );
  NAND2X0 U6137 ( .IN1(n3524), .IN2(n1470), .QN(n3551) );
  NAND2X0 U6138 ( .IN1(n3524), .IN2(n1464), .QN(n3642) );
  INVX0 U6139 ( .IN(n4815), .QN(n1421) );
  INVX0 U6140 ( .IN(n3312), .QN(n1788) );
  INVX0 U6141 ( .IN(n3315), .QN(n1794) );
  NAND2X0 U6142 ( .IN1(n1855), .IN2(n3623), .QN(n3625) );
  INVX0 U6143 ( .IN(n3314), .QN(n1795) );
  NAND2X0 U6144 ( .IN1(n1745), .IN2(n3549), .QN(n3552) );
  INVX0 U6145 ( .IN(n3470), .QN(n1437) );
  INVX0 U6146 ( .IN(n5102), .QN(n1448) );
  INVX0 U6147 ( .IN(n3550), .QN(n1470) );
  INVX0 U6148 ( .IN(n4361), .QN(n1440) );
  INVX0 U6149 ( .IN(n4209), .QN(n1430) );
  INVX0 U6150 ( .IN(n4270), .QN(n1434) );
  INVX0 U6151 ( .IN(n4255), .QN(n1433) );
  INVX0 U6152 ( .IN(n4225), .QN(n1431) );
  INVX0 U6153 ( .IN(n4331), .QN(n1438) );
  INVX0 U6154 ( .IN(n4346), .QN(n1439) );
  INVX0 U6155 ( .IN(n4240), .QN(n1432) );
  INVX0 U6156 ( .IN(n5120), .QN(n1443) );
  INVX0 U6157 ( .IN(n2712), .QN(n1411) );
  INVX0 U6158 ( .IN(n5110), .QN(n1442) );
  INVX0 U6159 ( .IN(n3003), .QN(n1464) );
  INVX0 U6160 ( .IN(n3007), .QN(n1471) );
  INVX0 U6161 ( .IN(n3337), .QN(n1800) );
  INVX0 U6162 ( .IN(n3569), .QN(n1469) );
  INVX0 U6163 ( .IN(n6027), .QN(n1402) );
  INVX0 U6164 ( .IN(n2723), .QN(n1474) );
  INVX0 U6165 ( .IN(n3606), .QN(n1467) );
  INVX0 U6166 ( .IN(n3588), .QN(n1468) );
  INVX0 U6167 ( .IN(n3165), .QN(n1482) );
  INVX0 U6168 ( .IN(n2398), .QN(n1802) );
  INVX0 U6169 ( .IN(n3352), .QN(n1791) );
  INVX0 U6170 ( .IN(n3311), .QN(n1790) );
  INVX0 U6171 ( .IN(n2449), .QN(n1423) );
  INVX0 U6172 ( .IN(n2545), .QN(n1801) );
  INVX0 U6173 ( .IN(n3208), .QN(n1367) );
  INVX0 U6174 ( .IN(n3107), .QN(n1335) );
  INVX0 U6175 ( .IN(n3127), .QN(n1327) );
  INVX0 U6176 ( .IN(n3148), .QN(n1319) );
  INVX0 U6177 ( .IN(n3188), .QN(n1376) );
  INVX0 U6178 ( .IN(n3228), .QN(n1358) );
  INVX0 U6179 ( .IN(n3167), .QN(n1311) );
  INVX0 U6180 ( .IN(n3246), .QN(n1349) );
  INVX0 U6181 ( .IN(n4541), .QN(n1441) );
  INVX0 U6182 ( .IN(n5233), .QN(n1446) );
  INVX0 U6183 ( .IN(n5211), .QN(n1444) );
  NAND2X0 U6184 ( .IN1(n1492), .IN2(n5962), .QN(n2416) );
  NAND2X0 U6185 ( .IN1(n1987), .IN2(n4194), .QN(n5087) );
  NAND2X0 U6186 ( .IN1(n3799), .IN2(n1843), .QN(n3503) );
  NAND2X0 U6187 ( .IN1(n2101), .IN2(n1558), .QN(n2676) );
  NAND2X0 U6188 ( .IN1(n2135), .IN2(n1704), .QN(n2655) );
  NAND2X0 U6189 ( .IN1(n2136), .IN2(n1704), .QN(n2659) );
  NAND2X0 U6190 ( .IN1(n2103), .IN2(n1558), .QN(n2680) );
  NAND2X0 U6191 ( .IN1(n3799), .IN2(n1842), .QN(n3474) );
  NAND2X0 U6192 ( .IN1(n3799), .IN2(n1845), .QN(n3484) );
  NAND2X0 U6193 ( .IN1(n3799), .IN2(n1844), .QN(n3399) );
  NAND2X0 U6194 ( .IN1(n1499), .IN2(g31863), .QN(n4159) );
  NAND2X0 U6195 ( .IN1(n1661), .IN2(n1770), .QN(n4133) );
  NAND2X0 U6196 ( .IN1(n2228), .IN2(n1859), .QN(n4121) );
  NAND2X0 U6197 ( .IN1(n2072), .IN2(n1762), .QN(n4085) );
  NAND2X0 U6198 ( .IN1(n1670), .IN2(n1713), .QN(n4073) );
  NAND2X0 U6199 ( .IN1(n2218), .IN2(n1499), .QN(n4157) );
  NAND2X0 U6200 ( .IN1(n2131), .IN2(n1863), .QN(n4109) );
  AND3X1 U6201 ( .IN1(n3033), .IN2(n1488), .IN3(n1565), .Q(n3024) );
  AND3X1 U6202 ( .IN1(n3033), .IN2(n1484), .IN3(n1611), .Q(n3066) );
  NOR2X0 U6203 ( .IN1(n3588), .IN2(n3592), .QN(n3591) );
  NOR2X0 U6204 ( .IN1(n3606), .IN2(n3610), .QN(n3609) );
  NOR2X0 U6205 ( .IN1(n3007), .IN2(n3535), .QN(n3534) );
  NOR2X0 U6206 ( .IN1(n3006), .IN2(n3516), .QN(n3515) );
  INVX0 U6207 ( .IN(n3592), .QN(n1859) );
  INVX0 U6208 ( .IN(n3516), .QN(n1713) );
  INVX0 U6209 ( .IN(n3610), .QN(n1770) );
  INVX0 U6210 ( .IN(n3535), .QN(n1762) );
  ISOLANDX1 U6211 ( .D(n3623), .ISO(n1466), .Q(n3622) );
  ISOLANDX1 U6212 ( .D(n3587), .ISO(n3588), .Q(n3586) );
  ISOLANDX1 U6213 ( .D(n3605), .ISO(n3606), .Q(n3604) );
  ISOLANDX1 U6214 ( .D(n3568), .ISO(n3569), .Q(n3567) );
  ISOLANDX1 U6215 ( .D(n3549), .ISO(n3550), .Q(n3548) );
  ISOLANDX1 U6216 ( .D(n3512), .ISO(n3006), .Q(n3511) );
  ISOLANDX1 U6217 ( .D(n3531), .ISO(n3007), .Q(n3530) );
  ISOLANDX1 U6218 ( .D(n3641), .ISO(n3003), .Q(n3640) );
  NOR2X0 U6219 ( .IN1(n3003), .IN2(n3645), .QN(n3644) );
  NOR2X0 U6220 ( .IN1(n3569), .IN2(n3573), .QN(n3572) );
  NOR2X0 U6221 ( .IN1(n2723), .IN2(n1599), .QN(n3244) );
  INVX0 U6222 ( .IN(n3645), .QN(n1499) );
  INVX0 U6223 ( .IN(n3573), .QN(n1863) );
  INVX0 U6224 ( .IN(n4333), .QN(n1502) );
  INVX0 U6225 ( .IN(n4227), .QN(n1566) );
  INVX0 U6226 ( .IN(n4272), .QN(n1559) );
  INVX0 U6227 ( .IN(n4363), .QN(n1589) );
  INVX0 U6228 ( .IN(n4257), .QN(n1561) );
  INVX0 U6229 ( .IN(n4212), .QN(n1674) );
  INVX0 U6230 ( .IN(n4242), .QN(n1563) );
  INVX0 U6231 ( .IN(n4348), .QN(n1594) );
  INVX0 U6232 ( .IN(n5063), .QN(n1574) );
  NAND2X0 U6233 ( .IN1(n1859), .IN2(n3587), .QN(n3590) );
  NAND2X0 U6234 ( .IN1(n1770), .IN2(n3605), .QN(n3608) );
  NAND2X0 U6235 ( .IN1(n1762), .IN2(n3531), .QN(n3533) );
  NAND2X0 U6236 ( .IN1(n1863), .IN2(n3568), .QN(n3571) );
  NAND2X0 U6237 ( .IN1(n1499), .IN2(n3641), .QN(n3643) );
  NAND2X0 U6238 ( .IN1(n1713), .IN2(n3512), .QN(n3514) );
  INVX0 U6239 ( .IN(n3286), .QN(n1844) );
  INVX0 U6240 ( .IN(n2579), .QN(n1298) );
  INVX0 U6241 ( .IN(n2755), .QN(n1306) );
  INVX0 U6242 ( .IN(n2770), .QN(n1302) );
  INVX0 U6243 ( .IN(n3439), .QN(n1284) );
  INVX0 U6244 ( .IN(n3429), .QN(n1285) );
  INVX0 U6245 ( .IN(n3419), .QN(n1286) );
  INVX0 U6246 ( .IN(n3409), .QN(n1287) );
  INVX0 U6247 ( .IN(n4687), .QN(n1883) );
  INVX0 U6248 ( .IN(n4658), .QN(n1890) );
  INVX0 U6249 ( .IN(n4612), .QN(n1866) );
  INVX0 U6250 ( .IN(n4635), .QN(n2305) );
  INVX0 U6251 ( .IN(n4677), .QN(n1748) );
  INVX0 U6252 ( .IN(n4566), .QN(n2119) );
  INVX0 U6253 ( .IN(n4682), .QN(n1943) );
  INVX0 U6254 ( .IN(n4589), .QN(n1621) );
  INVX0 U6255 ( .IN(n4801), .QN(n1571) );
  INVX0 U6256 ( .IN(n4050), .QN(n1864) );
  INVX0 U6257 ( .IN(n3242), .QN(n1289) );
  INVX0 U6258 ( .IN(n2735), .QN(n1486) );
  INVX0 U6259 ( .IN(n3162), .QN(n1293) );
  INVX0 U6260 ( .IN(n3183), .QN(n1292) );
  INVX0 U6261 ( .IN(n3223), .QN(n1290) );
  INVX0 U6262 ( .IN(n3143), .QN(n1294) );
  INVX0 U6263 ( .IN(n3203), .QN(n1291) );
  INVX0 U6264 ( .IN(n2738), .QN(n1487) );
  INVX0 U6265 ( .IN(n3005), .QN(n1466) );
  INVX0 U6266 ( .IN(n4808), .QN(n1986) );
  INVX0 U6267 ( .IN(n3131), .QN(n1295) );
  INVX0 U6268 ( .IN(n3111), .QN(n1296) );
  INVX0 U6269 ( .IN(n4176), .QN(n1837) );
  INVX0 U6270 ( .IN(n4194), .QN(n1927) );
  INVX0 U6271 ( .IN(n3907), .QN(n1577) );
  INVX0 U6272 ( .IN(n3773), .QN(n2225) );
  INVX0 U6273 ( .IN(n3807), .QN(n1510) );
  INVX0 U6274 ( .IN(n3950), .QN(n1904) );
  INVX0 U6275 ( .IN(n3841), .QN(n1817) );
  INVX0 U6276 ( .IN(n3983), .QN(n1681) );
  INVX0 U6277 ( .IN(n3874), .QN(n1969) );
  INVX0 U6278 ( .IN(n4014), .QN(n1731) );
  ISOLANDX1 U6279 ( .D(n4537), .ISO(n5337), .Q(n4201) );
  ISOLANDX1 U6280 ( .D(n4201), .ISO(n5336), .Q(n3745) );
  ISOLANDX1 U6281 ( .D(n3745), .ISO(n5294), .Q(n3684) );
  ISOLANDX1 U6282 ( .D(n3684), .ISO(n5552), .Q(n3274) );
  ISOLANDX1 U6283 ( .D(n3274), .ISO(n5472), .Q(n2982) );
  ISOLANDX1 U6284 ( .D(n2982), .ISO(n5476), .Q(n2706) );
  ISOLANDX1 U6285 ( .D(n2706), .ISO(n5550), .Q(n2649) );
  ISOLANDX1 U6286 ( .D(n2649), .ISO(n5473), .Q(n2556) );
  ISOLANDX1 U6287 ( .D(n2556), .ISO(n5475), .Q(n2509) );
  ISOLANDX1 U6288 ( .D(n2509), .ISO(n5474), .Q(n2487) );
  ISOLANDX1 U6289 ( .D(n2487), .ISO(n5339), .Q(n2427) );
  ISOLANDX1 U6290 ( .D(n2427), .ISO(n5672), .Q(n2423) );
  ISOLANDX1 U6291 ( .D(n4826), .ISO(n5335), .Q(n4537) );
  ISOLANDX1 U6292 ( .D(n4959), .ISO(n6145), .Q(n2421) );
  INVX0 U6293 ( .IN(n6683), .QN(n6679) );
  INVX0 U6294 ( .IN(n4872), .QN(n1648) );
  AO21X1 U6295 ( .IN1(n4172), .IN2(n2034), .IN3(n4173), .Q(n4169) );
  AO21X1 U6296 ( .IN1(n4190), .IN2(n1696), .IN3(n4191), .Q(n4187) );
  AND3X1 U6297 ( .IN1(n4894), .IN2(n4895), .IN3(n6024), .Q(n4172) );
  AND3X1 U6298 ( .IN1(n4919), .IN2(n4920), .IN3(n6021), .Q(n4190) );
  AO22X1 U6299 ( .IN1(n4871), .IN2(n6268), .IN3(n4864), .IN4(n4872), .Q(n4859)
         );
  OA21X1 U6300 ( .IN1(n4169), .IN2(n4171), .IN3(n6409), .Q(g30344) );
  XNOR2X1 U6301 ( .IN1(n5364), .IN2(n6024), .Q(n4171) );
  OA21X1 U6302 ( .IN1(n4187), .IN2(n4189), .IN3(n6410), .Q(g30338) );
  XNOR2X1 U6303 ( .IN1(n5363), .IN2(n6021), .Q(n4189) );
  OA21X1 U6304 ( .IN1(n2775), .IN2(n2761), .IN3(n2714), .Q(n2730) );
  NAND3X0 U6305 ( .IN1(n1700), .IN2(n2761), .IN3(n1609), .QN(n3010) );
  NAND3X0 U6306 ( .IN1(n1554), .IN2(n2775), .IN3(n1728), .QN(n3011) );
  NAND2X0 U6307 ( .IN1(n2730), .IN2(n2428), .QN(g34425) );
  AO21X1 U6308 ( .IN1(n4062), .IN2(n4455), .IN3(n4411), .Q(n3627) );
  NAND2X0 U6309 ( .IN1(n4388), .IN2(n5378), .QN(n4455) );
  AO21X1 U6310 ( .IN1(n4062), .IN2(n4410), .IN3(n4411), .Q(n3554) );
  NAND2X0 U6311 ( .IN1(n4388), .IN2(n5379), .QN(n4410) );
  NOR2X0 U6312 ( .IN1(n4845), .IN2(n4843), .QN(n4842) );
  NAND2X0 U6313 ( .IN1(n4838), .IN2(n4839), .QN(g28030) );
  NAND3X0 U6314 ( .IN1(n4850), .IN2(n1425), .IN3(n4842), .QN(n4838) );
  NAND4X0 U6315 ( .IN1(n4840), .IN2(n1426), .IN3(n1427), .IN4(n2469), .QN(
        n4839) );
  INVX0 U6316 ( .IN(n2471), .QN(n1425) );
  NAND2X0 U6317 ( .IN1(n3751), .IN2(n3752), .QN(g31793) );
  NAND4X0 U6318 ( .IN1(n2477), .IN2(n3762), .IN3(n2479), .IN4(n2474), .QN(
        n3751) );
  NAND4X0 U6319 ( .IN1(n3753), .IN2(n2478), .IN3(n2475), .IN4(n2473), .QN(
        n3752) );
  AO22X1 U6320 ( .IN1(n3763), .IN2(n2473), .IN3(n2478), .IN4(n2475), .Q(n3762)
         );
  AND3X1 U6321 ( .IN1(n1489), .IN2(n5323), .IN3(n3060), .Q(n2775) );
  NOR2X0 U6322 ( .IN1(g34977), .IN2(n6077), .QN(n2525) );
  OA222X1 U6323 ( .IN1(n3304), .IN2(n3305), .IN3(n3306), .IN4(n5483), .IN5(
        n3307), .IN6(n5341), .Q(n3303) );
  OA222X1 U6324 ( .IN1(n3304), .IN2(n3305), .IN3(n3306), .IN4(n5290), .IN5(
        n3307), .IN6(n5329), .Q(n3325) );
  OA221X1 U6325 ( .IN1(n3307), .IN2(n5478), .IN3(n3306), .IN4(n5343), .IN5(
        n3333), .Q(n3332) );
  OA221X1 U6326 ( .IN1(n3307), .IN2(n5328), .IN3(n3306), .IN4(n5289), .IN5(
        n3333), .Q(n3343) );
  INVX0 U6327 ( .IN(n6678), .QN(n6677) );
  INVX0 U6328 ( .IN(n6682), .QN(n6681) );
  INVX0 U6329 ( .IN(g34977), .QN(n1453) );
  INVX0 U6330 ( .IN(g34979), .QN(n1309) );
  AO22X1 U6331 ( .IN1(n2479), .IN2(n2477), .IN3(n2474), .IN4(n3754), .Q(n3753)
         );
  AO21X1 U6332 ( .IN1(n2479), .IN2(n3755), .IN3(n2477), .Q(n3754) );
  OAI21X1 U6333 ( .IN1(n1417), .IN2(n3756), .IN3(n3757), .QN(n3755) );
  AOI22X1 U6334 ( .IN1(n3758), .IN2(n3759), .IN3(n3760), .IN4(n3761), .QN(
        n3756) );
  INVX0 U6335 ( .IN(g34978), .QN(n1452) );
  AO22X1 U6336 ( .IN1(n4851), .IN2(n2469), .IN3(n1426), .IN4(n1427), .Q(n4850)
         );
  NAND2X0 U6337 ( .IN1(n4852), .IN2(n4853), .QN(n4851) );
  ISOLANDX1 U6338 ( .D(n4210), .ISO(n6144), .Q(n3765) );
  INVX0 U6339 ( .IN(g34971), .QN(n1277) );
  INVX0 U6340 ( .IN(g34975), .QN(n1455) );
  ISOLANDX1 U6341 ( .D(n6034), .ISO(n3479), .Q(n3951) );
  ISOLANDX1 U6342 ( .D(n6029), .ISO(n3404), .Q(n3774) );
  ISOLANDX1 U6343 ( .D(n6032), .ISO(n3424), .Q(n3842) );
  ISOLANDX1 U6344 ( .D(n6031), .ISO(n3414), .Q(n3808) );
  ISOLANDX1 U6345 ( .D(n6034), .ISO(n3444), .Q(n3908) );
  ISOLANDX1 U6346 ( .D(n6033), .ISO(n3489), .Q(n3984) );
  ISOLANDX1 U6347 ( .D(n6032), .ISO(n3434), .Q(n3875) );
  ISOLANDX1 U6348 ( .D(n6030), .ISO(n3500), .Q(n4015) );
  ISOLANDX1 U6349 ( .D(n6033), .ISO(n3446), .Q(n3914) );
  ISOLANDX1 U6350 ( .D(n6029), .ISO(n3406), .Q(n3780) );
  ISOLANDX1 U6351 ( .D(n6032), .ISO(n3481), .Q(n3957) );
  ISOLANDX1 U6352 ( .D(n6032), .ISO(n3426), .Q(n3848) );
  ISOLANDX1 U6353 ( .D(n6031), .ISO(n3491), .Q(n3990) );
  ISOLANDX1 U6354 ( .D(n6031), .ISO(n3416), .Q(n3814) );
  ISOLANDX1 U6355 ( .D(n6033), .ISO(n3436), .Q(n3881) );
  ISOLANDX1 U6356 ( .D(n6030), .ISO(n3502), .Q(n4022) );
  ISOLANDX1 U6357 ( .D(n6029), .ISO(n3501), .Q(n4027) );
  ISOLANDX1 U6358 ( .D(n6030), .ISO(n3407), .Q(n3785) );
  ISOLANDX1 U6359 ( .D(n6029), .ISO(n3482), .Q(n3962) );
  ISOLANDX1 U6360 ( .D(n6033), .ISO(n3427), .Q(n3853) );
  ISOLANDX1 U6361 ( .D(n6034), .ISO(n3437), .Q(n3886) );
  ISOLANDX1 U6362 ( .D(n6030), .ISO(n3417), .Q(n3819) );
  ISOLANDX1 U6363 ( .D(n6031), .ISO(n3492), .Q(n3995) );
  ISOLANDX1 U6364 ( .D(n6034), .ISO(n3447), .Q(n3919) );
  ISOLANDX1 U6365 ( .D(n3682), .ISO(n5471), .Q(n3272) );
  ISOLANDX1 U6366 ( .D(n3272), .ISO(n5331), .Q(n2980) );
  ISOLANDX1 U6367 ( .D(n2980), .ISO(n5332), .Q(n2704) );
  ISOLANDX1 U6368 ( .D(n2704), .ISO(n5333), .Q(n2647) );
  ISOLANDX1 U6369 ( .D(n2647), .ISO(n5334), .Q(n2554) );
  ISOLANDX1 U6370 ( .D(n2554), .ISO(n5330), .Q(n2507) );
  ISOLANDX1 U6371 ( .D(n2507), .ISO(n5551), .Q(n2485) );
  ISOLANDX1 U6372 ( .D(n2485), .ISO(n5293), .Q(n2425) );
  ISOLANDX1 U6373 ( .D(n2425), .ISO(n5292), .Q(n2419) );
  ISOLANDX1 U6374 ( .D(n3743), .ISO(n5470), .Q(n3682) );
  ISOLANDX1 U6375 ( .D(n2419), .ISO(n5291), .Q(n2405) );
  OR3X1 U6376 ( .IN1(n4848), .IN2(n4846), .IN3(n4849), .Q(n4845) );
  INVX0 U6377 ( .IN(g34970), .QN(n1457) );
  INVX0 U6378 ( .IN(g34974), .QN(n1456) );
  NAND3X0 U6379 ( .IN1(n3760), .IN2(n3758), .IN3(n3761), .QN(n3757) );
  INVX0 U6380 ( .IN(g34976), .QN(n1454) );
  INVX0 U6381 ( .IN(n4955), .QN(n1539) );
  OAI21X1 U6382 ( .IN1(n2471), .IN2(n4841), .IN3(n1424), .QN(n4840) );
  OA21X1 U6383 ( .IN1(n4843), .IN2(n4844), .IN3(n4845), .Q(n4841) );
  OA22X1 U6384 ( .IN1(n4846), .IN2(n4847), .IN3(n4848), .IN4(n4849), .Q(n4844)
         );
  AND2X1 U6385 ( .IN1(n4849), .IN2(n4848), .Q(n4847) );
  XNOR2X1 U6386 ( .IN1(g34977), .IN2(n1452), .Q(n2402) );
  XNOR2X1 U6387 ( .IN1(g34975), .IN2(n1454), .Q(n2403) );
  OR2X1 U6388 ( .IN1(n3761), .IN2(n3760), .Q(n3759) );
  INVX0 U6389 ( .IN(n4326), .QN(n2102) );
  INVX0 U6390 ( .IN(n4304), .QN(n2134) );
  INVX0 U6391 ( .IN(n2690), .QN(n1728) );
  INVX0 U6392 ( .IN(n2670), .QN(n1609) );
  INVX0 U6393 ( .IN(n2393), .QN(n1278) );
  INVX0 U6394 ( .IN(n5125), .QN(n2077) );
  INVX0 U6395 ( .IN(n3764), .QN(n1417) );
  NOR2X0 U6396 ( .IN1(n6082), .IN2(n2760), .QN(n3098) );
  AO21X1 U6397 ( .IN1(n4062), .IN2(n4433), .IN3(n4052), .Q(n3592) );
  NAND2X0 U6398 ( .IN1(n4388), .IN2(n5610), .QN(n4433) );
  AO21X1 U6399 ( .IN1(n4062), .IN2(n4387), .IN3(n4052), .Q(n3516) );
  NAND2X0 U6400 ( .IN1(n4388), .IN2(n5609), .QN(n4387) );
  NAND4X0 U6401 ( .IN1(n2715), .IN2(n2716), .IN3(n2717), .IN4(n2718), .QN(
        g34843) );
  NOR4X0 U6402 ( .IN1(n2719), .IN2(n2720), .IN3(n2721), .IN4(n2722), .QN(n2718) );
  OA21X1 U6403 ( .IN1(n2723), .IN2(n2724), .IN3(n2725), .Q(n2717) );
  NAND2X0 U6404 ( .IN1(n2760), .IN2(n6169), .QN(n2615) );
  NAND2X0 U6405 ( .IN1(n3392), .IN2(n3381), .QN(n3312) );
  NAND2X0 U6406 ( .IN1(n2531), .IN2(n2552), .QN(n3315) );
  NAND2X0 U6407 ( .IN1(n3391), .IN2(n2552), .QN(n3314) );
  NOR2X0 U6408 ( .IN1(n4946), .IN2(n6065), .QN(n4944) );
  NAND2X0 U6409 ( .IN1(n6221), .IN2(n3296), .QN(n4361) );
  NAND2X0 U6410 ( .IN1(n6184), .IN2(n3287), .QN(n4270) );
  NAND2X0 U6411 ( .IN1(n6209), .IN2(n3295), .QN(n4209) );
  NAND2X0 U6412 ( .IN1(n6202), .IN2(n3289), .QN(n4255) );
  NAND2X0 U6413 ( .IN1(n6206), .IN2(n3292), .QN(n4225) );
  NAND2X0 U6414 ( .IN1(n6235), .IN2(n3298), .QN(n4331) );
  NAND2X0 U6415 ( .IN1(n6231), .IN2(n3299), .QN(n4346) );
  NAND2X0 U6416 ( .IN1(n6207), .IN2(n3294), .QN(n4240) );
  ISOLANDX1 U6417 ( .D(n4198), .ISO(n6144), .Q(n2404) );
  NOR2X0 U6418 ( .IN1(n6081), .IN2(g28753), .QN(n3057) );
  NAND2X0 U6419 ( .IN1(n6668), .IN2(n4821), .QN(n4815) );
  AND3X1 U6420 ( .IN1(n4890), .IN2(n2631), .IN3(n4888), .Q(n4889) );
  NAND2X0 U6421 ( .IN1(n5300), .IN2(n5516), .QN(n4890) );
  NAND3X0 U6422 ( .IN1(n5299), .IN2(n5465), .IN3(n4466), .QN(n3645) );
  AO21X1 U6423 ( .IN1(n4388), .IN2(n5544), .IN3(n2048), .Q(n4466) );
  OA21X1 U6424 ( .IN1(n2962), .IN2(n5526), .IN3(n2963), .Q(n2956) );
  OA21X1 U6425 ( .IN1(n5526), .IN2(n2916), .IN3(n2917), .Q(n2910) );
  OA21X1 U6426 ( .IN1(n5757), .IN2(n2822), .IN3(n2823), .Q(n2816) );
  OA21X1 U6427 ( .IN1(n2868), .IN2(n5757), .IN3(n2869), .Q(n2862) );
  NAND3X0 U6428 ( .IN1(n5299), .IN2(n5465), .IN3(n4422), .QN(n3573) );
  AO21X1 U6429 ( .IN1(n4388), .IN2(n5545), .IN3(n2048), .Q(n4422) );
  NAND2X0 U6430 ( .IN1(n3653), .IN2(n3581), .QN(n3003) );
  AND3X1 U6431 ( .IN1(n3381), .IN2(n5324), .IN3(n3382), .Q(n2459) );
  NAND2X0 U6432 ( .IN1(n2439), .IN2(n2440), .QN(g26876) );
  NAND2X0 U6433 ( .IN1(n2432), .IN2(n2433), .QN(g26877) );
  NAND2X0 U6434 ( .IN1(n1423), .IN2(n2447), .QN(g28042) );
  NAND3X0 U6435 ( .IN1(n3381), .IN2(n5468), .IN3(n2531), .QN(n3311) );
  NAND2X0 U6436 ( .IN1(n6214), .IN2(n5729), .QN(n3470) );
  NAND2X0 U6437 ( .IN1(n3543), .IN2(n3525), .QN(n3007) );
  AND3X1 U6438 ( .IN1(n5324), .IN2(n5469), .IN3(n3396), .Q(n2531) );
  NAND2X0 U6439 ( .IN1(n6191), .IN2(n4824), .QN(n5120) );
  NAND2X0 U6440 ( .IN1(n6212), .IN2(n4499), .QN(n5233) );
  NAND3X0 U6441 ( .IN1(n3381), .IN2(n5468), .IN3(n2528), .QN(n3352) );
  NAND2X0 U6442 ( .IN1(n3562), .IN2(n3525), .QN(n3550) );
  NAND2X0 U6443 ( .IN1(n6192), .IN2(n4818), .QN(n5110) );
  NAND2X0 U6444 ( .IN1(n6193), .IN2(n4475), .QN(n5211) );
  NAND2X0 U6445 ( .IN1(n5948), .IN2(n6025), .QN(n3321) );
  ISOLANDX1 U6446 ( .D(n6022), .ISO(n1300), .Q(n3524) );
  NAND2X0 U6447 ( .IN1(n3750), .IN2(n6167), .QN(n2712) );
  NOR2X0 U6448 ( .IN1(n5524), .IN2(n2800), .QN(n2806) );
  NOR2X0 U6449 ( .IN1(n5523), .IN2(n2824), .QN(n2830) );
  NOR2X0 U6450 ( .IN1(n5513), .IN2(n2847), .QN(n2853) );
  NOR2X0 U6451 ( .IN1(n5514), .IN2(n2870), .QN(n2876) );
  NAND2X0 U6452 ( .IN1(n2761), .IN2(n5298), .QN(n2735) );
  NAND2X0 U6453 ( .IN1(n4962), .IN2(n6157), .QN(n4541) );
  NAND2X0 U6454 ( .IN1(n2775), .IN2(n5298), .QN(n2738) );
  NAND2X0 U6455 ( .IN1(n4948), .IN2(n6165), .QN(n5102) );
  NOR2X0 U6456 ( .IN1(n2669), .IN2(n6063), .QN(n2759) );
  NAND3X0 U6457 ( .IN1(n5356), .IN2(n5538), .IN3(n1313), .QN(n3167) );
  NAND3X0 U6458 ( .IN1(n5351), .IN2(n5521), .IN3(n1337), .QN(n3107) );
  NAND3X0 U6459 ( .IN1(n5357), .IN2(n5522), .IN3(n1329), .QN(n3127) );
  NAND3X0 U6460 ( .IN1(n5353), .IN2(n5537), .IN3(n1321), .QN(n3148) );
  NAND3X0 U6461 ( .IN1(n5354), .IN2(n5534), .IN3(n2930), .QN(n3208) );
  NAND3X0 U6462 ( .IN1(n5352), .IN2(n5536), .IN3(n2953), .QN(n3228) );
  NAND3X0 U6463 ( .IN1(n5355), .IN2(n5535), .IN3(n2906), .QN(n3188) );
  NAND3X0 U6464 ( .IN1(n5362), .IN2(n5598), .IN3(n2966), .QN(n3246) );
  ISOLANDX1 U6465 ( .D(n3653), .ISO(n5600), .Q(n4388) );
  NAND2X0 U6466 ( .IN1(n6680), .IN2(n5630), .QN(n2449) );
  NAND2X0 U6467 ( .IN1(n3394), .IN2(n3392), .QN(n2545) );
  NOR2X0 U6468 ( .IN1(n2592), .IN2(n6078), .QN(n2591) );
  NOR2X0 U6469 ( .IN1(n5538), .IN2(n2870), .QN(n2873) );
  NOR2X0 U6470 ( .IN1(n5521), .IN2(n2800), .QN(n2803) );
  NOR2X0 U6471 ( .IN1(n5522), .IN2(n2824), .QN(n2827) );
  NOR2X0 U6472 ( .IN1(n5537), .IN2(n2847), .QN(n2850) );
  NAND3X0 U6473 ( .IN1(n2713), .IN2(n1475), .IN3(n2714), .QN(g34383) );
  NAND4X0 U6474 ( .IN1(n2726), .IN2(n2727), .IN3(n2728), .IN4(n2729), .QN(
        n2713) );
  INVX0 U6475 ( .IN(g34843), .QN(n1475) );
  NOR2X0 U6476 ( .IN1(n1482), .IN2(n1483), .QN(n2728) );
  NAND3X0 U6477 ( .IN1(n2993), .IN2(n1465), .IN3(n2714), .QN(g34201) );
  NAND4X0 U6478 ( .IN1(n3006), .IN2(n3007), .IN3(n3008), .IN4(n3009), .QN(
        n2993) );
  INVX0 U6479 ( .IN(g34781), .QN(n1465) );
  NOR4X0 U6480 ( .IN1(n1464), .IN2(n3005), .IN3(n1467), .IN4(n1468), .QN(n3009) );
  OAI22X1 U6481 ( .IN1(n6306), .IN2(n5787), .IN3(n2801), .IN4(n6142), .QN(
        g34019) );
  OA22X1 U6482 ( .IN1(n2792), .IN2(n2802), .IN3(n1341), .IN4(n5800), .Q(n2801)
         );
  INVX0 U6483 ( .IN(n2802), .QN(n1341) );
  NAND2X0 U6484 ( .IN1(n2803), .IN2(n5524), .QN(n2802) );
  NAND3X0 U6485 ( .IN1(n5519), .IN2(n5287), .IN3(n3195), .QN(n2723) );
  AND3X1 U6486 ( .IN1(n5516), .IN2(n5300), .IN3(n5349), .Q(n3653) );
  NAND3X0 U6487 ( .IN1(n3581), .IN2(n5300), .IN3(n3505), .QN(n3588) );
  NAND3X0 U6488 ( .IN1(n5349), .IN2(n5516), .IN3(n3525), .QN(n3569) );
  NAND3X0 U6489 ( .IN1(n3581), .IN2(n5300), .IN3(n3543), .QN(n3606) );
  NOR2X0 U6490 ( .IN1(n2689), .IN2(n6063), .QN(n2774) );
  NAND2X0 U6491 ( .IN1(n2548), .IN2(n1461), .QN(n3320) );
  AND2X1 U6492 ( .IN1(n3397), .IN2(n2531), .Q(n2548) );
  NAND2X0 U6493 ( .IN1(n2547), .IN2(n1461), .QN(n3317) );
  AND2X1 U6494 ( .IN1(n3397), .IN2(n3391), .Q(n2547) );
  AO21X1 U6495 ( .IN1(n6018), .IN2(n1492), .IN3(n6028), .Q(n3454) );
  AO21X1 U6496 ( .IN1(n6016), .IN2(n5962), .IN3(n6028), .Q(n3458) );
  ISOLANDX1 U6497 ( .D(n3581), .ISO(n3635), .Q(n3005) );
  NAND3X0 U6498 ( .IN1(n3382), .IN2(n5324), .IN3(n3394), .QN(n2398) );
  NOR2X0 U6499 ( .IN1(n6080), .IN2(n3079), .QN(n3081) );
  NOR2X0 U6500 ( .IN1(n6082), .IN2(n3018), .QN(n3020) );
  NOR2X0 U6501 ( .IN1(n6080), .IN2(n3088), .QN(n3091) );
  NOR2X0 U6502 ( .IN1(n6081), .IN2(n3047), .QN(n3049) );
  NOR2X0 U6503 ( .IN1(n6081), .IN2(n3038), .QN(n3040) );
  NAND3X0 U6504 ( .IN1(n2528), .IN2(n5468), .IN3(n3394), .QN(n3337) );
  OA21X1 U6505 ( .IN1(n4984), .IN2(n4985), .IN3(n6356), .Q(n2439) );
  NAND4X0 U6506 ( .IN1(n5410), .IN2(n5624), .IN3(n5279), .IN4(n5314), .QN(
        n4985) );
  NAND4X0 U6507 ( .IN1(n5411), .IN2(n5625), .IN3(n5278), .IN4(n5313), .QN(
        n4984) );
  NOR2X0 U6508 ( .IN1(n3069), .IN2(n6068), .QN(n3074) );
  NOR2X0 U6509 ( .IN1(n3027), .IN2(n6069), .QN(n3032) );
  OA21X1 U6510 ( .IN1(n4980), .IN2(n4981), .IN3(n6361), .Q(n2432) );
  NAND4X0 U6511 ( .IN1(n5620), .IN2(n5406), .IN3(n5310), .IN4(n5276), .QN(
        n4981) );
  NAND4X0 U6512 ( .IN1(n5619), .IN2(n5405), .IN3(n5311), .IN4(n5277), .QN(
        n4980) );
  OA222X1 U6513 ( .IN1(n3312), .IN2(n5334), .IN3(n3314), .IN4(n5472), .IN5(
        n3315), .IN6(n5288), .Q(n3327) );
  OA222X1 U6514 ( .IN1(n3352), .IN2(n5293), .IN3(n3314), .IN4(n5335), .IN5(
        n3315), .IN6(n5473), .Q(n3383) );
  OA222X1 U6515 ( .IN1(n3352), .IN2(n5291), .IN3(n3314), .IN4(n5336), .IN5(
        n3315), .IN6(n5474), .Q(n3359) );
  AND4X1 U6516 ( .IN1(n5323), .IN2(n5506), .IN3(n6418), .IN4(n5167), .Q(n5164)
         );
  AND3X1 U6517 ( .IN1(n5540), .IN2(n5348), .IN3(n5298), .Q(n5167) );
  NOR2X0 U6518 ( .IN1(n5549), .IN2(n1347), .QN(n2969) );
  NOR2X0 U6519 ( .IN1(n5516), .IN2(n5349), .QN(n3505) );
  NOR2X0 U6520 ( .IN1(n5362), .IN2(n1347), .QN(n2972) );
  NOR2X0 U6521 ( .IN1(n6080), .IN2(n3177), .QN(n2453) );
  NAND3X0 U6522 ( .IN1(n5519), .IN2(n5287), .IN3(n3116), .QN(n3165) );
  ISOLANDX1 U6523 ( .D(n4946), .ISO(n6145), .Q(n4945) );
  NOR2X0 U6524 ( .IN1(n6081), .IN2(n3254), .QN(n2455) );
  INVX0 U6525 ( .IN(n6683), .QN(n6680) );
  INVX0 U6526 ( .IN(n6678), .QN(n6676) );
  OA221X1 U6527 ( .IN1(n3311), .IN2(n5486), .IN3(n3312), .IN4(n5332), .IN5(
        n3351), .Q(n3346) );
  OA222X1 U6528 ( .IN1(n3352), .IN2(n5479), .IN3(n3314), .IN4(n5294), .IN5(
        n3315), .IN6(n5339), .Q(n3351) );
  NOR2X0 U6529 ( .IN1(n4527), .IN2(n6069), .QN(n4525) );
  NOR2X0 U6530 ( .IN1(n6083), .IN2(n4520), .QN(n4518) );
  OA221X1 U6531 ( .IN1(n5103), .IN2(n5104), .IN3(n5732), .IN4(n5105), .IN5(
        n6221), .Q(g25616) );
  NAND2X0 U6532 ( .IN1(n5104), .IN2(n4955), .QN(n5105) );
  NOR2X0 U6533 ( .IN1(n1539), .IN2(n5732), .QN(n5103) );
  XNOR3X1 U6534 ( .IN1(n5106), .IN2(n5107), .IN3(n5597), .Q(n5104) );
  NOR2X0 U6535 ( .IN1(n5380), .IN2(n2978), .QN(n2907) );
  NOR2X0 U6536 ( .IN1(n5535), .IN2(n1374), .QN(n2896) );
  NOR2X0 U6537 ( .IN1(n5536), .IN2(n1356), .QN(n2943) );
  NOR2X0 U6538 ( .IN1(n5534), .IN2(n1365), .QN(n2920) );
  AND3X1 U6539 ( .IN1(n1279), .IN2(n5652), .IN3(n5366), .Q(g30393) );
  AND3X1 U6540 ( .IN1(n5126), .IN2(n4835), .IN3(n6415), .Q(g25594) );
  NAND2X0 U6541 ( .IN1(n5627), .IN2(n4834), .QN(n5126) );
  ISOLANDX1 U6542 ( .D(n3581), .ISO(n5300), .Q(n3525) );
  NOR2X0 U6543 ( .IN1(n4821), .IN2(n6067), .QN(n4816) );
  NAND3X0 U6544 ( .IN1(n2528), .IN2(n1461), .IN3(n2552), .QN(n3345) );
  NAND3X0 U6545 ( .IN1(n2528), .IN2(n1461), .IN3(n2527), .QN(n3319) );
  NOR2X0 U6546 ( .IN1(n5282), .IN2(n6064), .QN(n4973) );
  NOR2X0 U6547 ( .IN1(n5321), .IN2(n6079), .QN(n4939) );
  NOR2X0 U6548 ( .IN1(n5322), .IN2(n6079), .QN(n4914) );
  NOR2X0 U6549 ( .IN1(n5710), .IN2(n6067), .QN(n4864) );
  NAND2X0 U6550 ( .IN1(n2550), .IN2(n1461), .QN(n3344) );
  AND3X1 U6551 ( .IN1(n2531), .IN2(n5468), .IN3(n3394), .Q(n2550) );
  ISOLANDX1 U6552 ( .D(n3281), .ISO(n5676), .Q(n3277) );
  ISOLANDX1 U6553 ( .D(n3276), .ISO(n5680), .Q(n2989) );
  ISOLANDX1 U6554 ( .D(n3277), .ISO(n5677), .Q(n2991) );
  ISOLANDX1 U6555 ( .D(n3687), .ISO(n5561), .Q(n3281) );
  ISOLANDX1 U6556 ( .D(n3279), .ISO(n5679), .Q(n3276) );
  NOR2X0 U6557 ( .IN1(n5964), .IN2(n6145), .QN(n2441) );
  AND4X1 U6558 ( .IN1(n5414), .IN2(n5631), .IN3(n5281), .IN4(n5316), .Q(n5964)
         );
  ISOLANDX1 U6559 ( .D(n2991), .ISO(n5678), .Q(n2710) );
  ISOLANDX1 U6560 ( .D(n2989), .ISO(n5675), .Q(n2707) );
  ISOLANDX1 U6561 ( .D(n3174), .ISO(n5327), .Q(n3116) );
  NAND4X0 U6562 ( .IN1(n2473), .IN2(n2474), .IN3(n2475), .IN4(n2476), .QN(
        n2437) );
  AND3X1 U6563 ( .IN1(n2477), .IN2(n2478), .IN3(n2479), .Q(n2476) );
  NAND4X0 U6564 ( .IN1(n1427), .IN2(n2469), .IN3(n1426), .IN4(n2470), .QN(
        n2438) );
  NOR2X0 U6565 ( .IN1(n2471), .IN2(n1424), .QN(n2470) );
  INVX0 U6566 ( .IN(n3269), .QN(n1447) );
  INVX0 U6567 ( .IN(n3261), .QN(n1445) );
  NOR2X0 U6568 ( .IN1(n4492), .IN2(n4495), .QN(n4494) );
  NOR2X0 U6569 ( .IN1(n4468), .IN2(n4471), .QN(n4470) );
  ISOLANDX1 U6570 ( .D(n3362), .ISO(n5477), .Q(n2527) );
  NAND3X0 U6571 ( .IN1(n3474), .IN2(n5648), .IN3(n6326), .QN(n3476) );
  NAND3X0 U6572 ( .IN1(n3399), .IN2(n5646), .IN3(n6326), .QN(n3401) );
  NAND3X0 U6573 ( .IN1(n3419), .IN2(n5649), .IN3(n6324), .QN(n3421) );
  NAND3X0 U6574 ( .IN1(n3429), .IN2(n5647), .IN3(n6325), .QN(n3431) );
  NAND3X0 U6575 ( .IN1(n3484), .IN2(n5645), .IN3(n6324), .QN(n3486) );
  NAND3X0 U6576 ( .IN1(n3439), .IN2(n5650), .IN3(n6326), .QN(n3441) );
  NAND3X0 U6577 ( .IN1(n3409), .IN2(n5651), .IN3(n6325), .QN(n3411) );
  NAND2X0 U6578 ( .IN1(n2546), .IN2(n1461), .QN(n3363) );
  NOR2X0 U6579 ( .IN1(n4824), .IN2(n6077), .QN(n5119) );
  NOR2X0 U6580 ( .IN1(n2618), .IN2(n6079), .QN(n2616) );
  NOR2X0 U6581 ( .IN1(n5390), .IN2(n6079), .QN(g25648) );
  OA21X1 U6582 ( .IN1(n2822), .IN2(n5755), .IN3(n2823), .Q(n2821) );
  OA21X1 U6583 ( .IN1(n5755), .IN2(n2868), .IN3(n2869), .Q(n2867) );
  OA21X1 U6584 ( .IN1(n2916), .IN2(n5756), .IN3(n2917), .Q(n2915) );
  OA21X1 U6585 ( .IN1(n5756), .IN2(n2962), .IN3(n2963), .Q(n2961) );
  NOR2X0 U6586 ( .IN1(n5568), .IN2(n6064), .QN(g25742) );
  NOR2X0 U6587 ( .IN1(n5563), .IN2(n6064), .QN(g25756) );
  NOR2X0 U6588 ( .IN1(n5569), .IN2(n6078), .QN(g25662) );
  NOR2X0 U6589 ( .IN1(n5567), .IN2(n6063), .QN(g25700) );
  NOR2X0 U6590 ( .IN1(n5566), .IN2(n6063), .QN(g25714) );
  NOR2X0 U6591 ( .IN1(n5564), .IN2(n6077), .QN(g25676) );
  NOR2X0 U6592 ( .IN1(n5565), .IN2(n6063), .QN(g25728) );
  NAND2X0 U6593 ( .IN1(n2536), .IN2(n1461), .QN(n3364) );
  AND2X1 U6594 ( .IN1(n3397), .IN2(n2528), .Q(n2536) );
  OA22X1 U6595 ( .IN1(n2738), .IN2(n2745), .IN3(n2740), .IN4(n2746), .Q(n2744)
         );
  OAI22X1 U6596 ( .IN1(n6316), .IN2(n5792), .IN3(n2964), .IN4(n6143), .QN(
        g33970) );
  OA22X1 U6597 ( .IN1(n2956), .IN2(n2965), .IN3(n1350), .IN4(n5791), .Q(n2964)
         );
  INVX0 U6598 ( .IN(n2965), .QN(n1350) );
  NAND2X0 U6599 ( .IN1(g31862), .IN2(n2966), .QN(n2965) );
  NBUFFX2 U6600 ( .IN(n3456), .Q(n6028) );
  OA22X1 U6601 ( .IN1(n5734), .IN2(n4268), .IN3(n4269), .IN4(n6048), .Q(g29285) );
  NAND2X0 U6602 ( .IN1(n4210), .IN2(n3287), .QN(n4268) );
  NOR2X0 U6603 ( .IN1(n4270), .IN2(n5734), .QN(n4269) );
  NBUFFX2 U6604 ( .IN(n3309), .Q(n6026) );
  NOR2X0 U6605 ( .IN1(n4475), .IN2(n4478), .QN(n4477) );
  OAI222X1 U6606 ( .IN1(n4543), .IN2(n5358), .IN3(n1715), .IN4(n4544), .IN5(
        n4545), .IN6(n5629), .QN(g29222) );
  INVX0 U6607 ( .IN(n3676), .QN(n1715) );
  NAND2X0 U6608 ( .IN1(n1448), .IN2(n5358), .QN(n4544) );
  OA21X1 U6609 ( .IN1(n3676), .IN2(n2076), .IN3(n6359), .Q(n4543) );
  OAI222X1 U6610 ( .IN1(n5517), .IN2(n2748), .IN3(n1307), .IN4(n2749), .IN5(
        n6300), .IN6(n5360), .QN(g34040) );
  OA22X1 U6611 ( .IN1(n2750), .IN2(n2751), .IN3(n6117), .IN4(n2752), .Q(n2749)
         );
  OAI222X1 U6612 ( .IN1(n5518), .IN2(n2763), .IN3(n1303), .IN4(n2764), .IN5(
        n6299), .IN6(n5361), .QN(g34032) );
  OA22X1 U6613 ( .IN1(n2765), .IN2(n2766), .IN3(n6117), .IN4(n2767), .Q(n2764)
         );
  OAI222X1 U6614 ( .IN1(n3501), .IN2(n1280), .IN3(n3502), .IN4(n3498), .IN5(
        n5366), .IN6(n6419), .QN(g33021) );
  INVX0 U6615 ( .IN(n4062), .QN(n2048) );
  NOR2X0 U6616 ( .IN1(n2759), .IN2(n5318), .QN(g34035) );
  NOR2X0 U6617 ( .IN1(n2759), .IN2(n5713), .QN(g34034) );
  NOR2X0 U6618 ( .IN1(n2759), .IN2(n5443), .QN(g34036) );
  NOR2X0 U6619 ( .IN1(n3674), .IN2(n6070), .QN(g32980) );
  OA22X1 U6620 ( .IN1(n1726), .IN2(n5754), .IN3(n2644), .IN4(n2645), .Q(n3674)
         );
  INVX0 U6621 ( .IN(n2645), .QN(n1726) );
  NOR2X0 U6622 ( .IN1(n6240), .IN2(n5750), .QN(g18597) );
  NOR2X0 U6623 ( .IN1(n6241), .IN2(n5710), .QN(g24298) );
  NOR2X0 U6624 ( .IN1(n2774), .IN2(n5440), .QN(g34027) );
  NOR2X0 U6625 ( .IN1(n2774), .IN2(n5712), .QN(g34026) );
  OAI21X1 U6626 ( .IN1(n5244), .IN2(n5562), .IN3(n6417), .QN(n5248) );
  NBUFFX2 U6627 ( .IN(n3456), .Q(n6027) );
  NAND2X0 U6628 ( .IN1(n3562), .IN2(n5300), .QN(n3635) );
  NOR2X0 U6629 ( .IN1(n3670), .IN2(n5731), .QN(g32982) );
  OA21X1 U6630 ( .IN1(n3254), .IN2(n3270), .IN3(n6405), .Q(n3670) );
  NOR2X0 U6631 ( .IN1(n3661), .IN2(n5730), .QN(g32985) );
  OA21X1 U6632 ( .IN1(n3177), .IN2(n3262), .IN3(n6406), .Q(n3661) );
  NBUFFX2 U6633 ( .IN(n3309), .Q(n6025) );
  OAI21X1 U6634 ( .IN1(n4818), .IN2(n4962), .IN3(n6418), .QN(n5116) );
  OR2X1 U6635 ( .IN1(n2475), .IN2(n2478), .Q(n3763) );
  OAI22X1 U6636 ( .IN1(n6316), .IN2(n5397), .IN3(n3043), .IN4(n3044), .QN(
        g33621) );
  OA22X1 U6637 ( .IN1(n3045), .IN2(n6119), .IN3(n1562), .IN4(n3046), .Q(n3044)
         );
  OA21X1 U6638 ( .IN1(n3047), .IN2(n5593), .IN3(n3048), .Q(n3045) );
  OAI22X1 U6639 ( .IN1(n6317), .IN2(n5398), .IN3(n3014), .IN4(n3015), .QN(
        g33627) );
  OA22X1 U6640 ( .IN1(n3016), .IN2(n6119), .IN3(n1705), .IN4(n3017), .Q(n3015)
         );
  OA21X1 U6641 ( .IN1(n3018), .IN2(n5590), .IN3(n3019), .Q(n3016) );
  OAI22X1 U6642 ( .IN1(n6314), .IN2(n5399), .IN3(n3075), .IN4(n3076), .QN(
        g33612) );
  OA22X1 U6643 ( .IN1(n3077), .IN2(n6119), .IN3(n1650), .IN4(n3078), .Q(n3076)
         );
  OA21X1 U6644 ( .IN1(n3079), .IN2(n5591), .IN3(n3080), .Q(n3077) );
  OAI22X1 U6645 ( .IN1(n6315), .IN2(n5395), .IN3(n3066), .IN4(n3067), .QN(
        g33614) );
  OA22X1 U6646 ( .IN1(n3068), .IN2(n6119), .IN3(n3069), .IN4(n3070), .Q(n3067)
         );
  OA21X1 U6647 ( .IN1(n1611), .IN2(n5594), .IN3(n3071), .Q(n3068) );
  OAI22X1 U6648 ( .IN1(n6316), .IN2(n5393), .IN3(n3052), .IN4(n3053), .QN(
        g33619) );
  OA22X1 U6649 ( .IN1(n3054), .IN2(n6119), .IN3(n1560), .IN4(n3055), .Q(n3053)
         );
  OA21X1 U6650 ( .IN1(g28753), .IN2(n5588), .IN3(n3056), .Q(n3054) );
  OAI22X1 U6651 ( .IN1(n6317), .IN2(n5394), .IN3(n3034), .IN4(n3035), .QN(
        g33623) );
  OA22X1 U6652 ( .IN1(n3036), .IN2(n6119), .IN3(n1564), .IN4(n3037), .Q(n3035)
         );
  OA21X1 U6653 ( .IN1(n3038), .IN2(n5589), .IN3(n3039), .Q(n3036) );
  OAI22X1 U6654 ( .IN1(n6317), .IN2(n5396), .IN3(n3024), .IN4(n3025), .QN(
        g33625) );
  OA22X1 U6655 ( .IN1(n3026), .IN2(n6119), .IN3(n3027), .IN4(n3028), .Q(n3025)
         );
  OA21X1 U6656 ( .IN1(n1565), .IN2(n5592), .IN3(n3029), .Q(n3026) );
  OAI22X1 U6657 ( .IN1(n6322), .IN2(n5343), .IN3(n4479), .IN4(n6141), .QN(
        g29237) );
  OA22X1 U6658 ( .IN1(n4480), .IN2(n4481), .IN3(n4482), .IN4(n5693), .Q(n4479)
         );
  NAND2X0 U6659 ( .IN1(n4472), .IN2(n4483), .QN(n4481) );
  NOR2X0 U6660 ( .IN1(n4480), .IN2(n4483), .QN(n4482) );
  OAI22X1 U6661 ( .IN1(n6323), .IN2(n5478), .IN3(n4503), .IN4(n6141), .QN(
        g29232) );
  OA22X1 U6662 ( .IN1(n4504), .IN2(n4505), .IN3(n4506), .IN4(n5692), .Q(n4503)
         );
  NAND2X0 U6663 ( .IN1(n4496), .IN2(n4507), .QN(n4505) );
  NOR2X0 U6664 ( .IN1(n4504), .IN2(n4507), .QN(n4506) );
  OAI22X1 U6665 ( .IN1(n4065), .IN2(n6146), .IN3(n4066), .IN4(n5777), .QN(
        g30387) );
  OA22X1 U6666 ( .IN1(n4067), .IN2(n4068), .IN3(n1712), .IN4(n5313), .Q(n4065)
         );
  OA21X1 U6667 ( .IN1(n5457), .IN2(n4067), .IN3(n6404), .Q(n4066) );
  NAND2X0 U6668 ( .IN1(n5457), .IN2(n5777), .QN(n4068) );
  OAI22X1 U6669 ( .IN1(n4101), .IN2(n6146), .IN3(n4102), .IN4(n5778), .QN(
        g30372) );
  OA22X1 U6670 ( .IN1(n4103), .IN2(n4104), .IN3(n1860), .IN4(n5624), .Q(n4101)
         );
  OA21X1 U6671 ( .IN1(n5458), .IN2(n4103), .IN3(n6406), .Q(n4102) );
  NAND2X0 U6672 ( .IN1(n5458), .IN2(n5778), .QN(n4104) );
  OAI22X1 U6673 ( .IN1(n4089), .IN2(n6146), .IN3(n4090), .IN4(n5779), .QN(
        g30377) );
  OA21X1 U6674 ( .IN1(n5459), .IN2(n4091), .IN3(n6405), .Q(n4090) );
  OA22X1 U6675 ( .IN1(n4091), .IN2(n4092), .IN3(n1742), .IN4(n5314), .Q(n4089)
         );
  NAND2X0 U6676 ( .IN1(n5459), .IN2(n5779), .QN(n4092) );
  OAI22X1 U6677 ( .IN1(n6320), .IN2(n5542), .IN3(n5210), .IN4(n6140), .QN(
        g24252) );
  OA22X1 U6678 ( .IN1(n5381), .IN2(n5302), .IN3(n6024), .IN4(n5577), .Q(n5210)
         );
  OAI22X1 U6679 ( .IN1(n6321), .IN2(n5329), .IN3(n4498), .IN4(n6141), .QN(
        g29233) );
  OA22X1 U6680 ( .IN1(n4499), .IN2(n4500), .IN3(n4501), .IN4(n5691), .Q(n4498)
         );
  NAND2X0 U6681 ( .IN1(n4496), .IN2(n4502), .QN(n4500) );
  NOR2X0 U6682 ( .IN1(n4499), .IN2(n4502), .QN(n4501) );
  OAI22X1 U6683 ( .IN1(n6303), .IN2(n5570), .IN3(n1284), .IN4(n3445), .QN(
        g33047) );
  OA21X1 U6684 ( .IN1(n6116), .IN2(n3446), .IN3(n3447), .Q(n3445) );
  OAI22X1 U6685 ( .IN1(n6305), .IN2(n5575), .IN3(n1285), .IN4(n3435), .QN(
        g33052) );
  OA21X1 U6686 ( .IN1(n6116), .IN2(n3436), .IN3(n3437), .Q(n3435) );
  OAI22X1 U6687 ( .IN1(n6302), .IN2(n5572), .IN3(n1282), .IN4(n3480), .QN(
        g33031) );
  OA21X1 U6688 ( .IN1(n6116), .IN2(n3481), .IN3(n3482), .Q(n3480) );
  OAI22X1 U6689 ( .IN1(n6305), .IN2(n5573), .IN3(n1286), .IN4(n3425), .QN(
        g33057) );
  OA21X1 U6690 ( .IN1(n6116), .IN2(n3426), .IN3(n3427), .Q(n3425) );
  OAI22X1 U6691 ( .IN1(n6306), .IN2(n5574), .IN3(n1287), .IN4(n3415), .QN(
        g33062) );
  OA21X1 U6692 ( .IN1(n6116), .IN2(n3416), .IN3(n3417), .Q(n3415) );
  OAI22X1 U6693 ( .IN1(n6306), .IN2(n5571), .IN3(n1283), .IN4(n3405), .QN(
        g33067) );
  OA21X1 U6694 ( .IN1(n6116), .IN2(n3406), .IN3(n3407), .Q(n3405) );
  OAI22X1 U6695 ( .IN1(n6301), .IN2(n5576), .IN3(n1281), .IN4(n3490), .QN(
        g33026) );
  OA21X1 U6696 ( .IN1(n6116), .IN2(n3491), .IN3(n3492), .Q(n3490) );
  OAI22X1 U6697 ( .IN1(n4149), .IN2(n6145), .IN3(n4150), .IN4(n5780), .QN(
        g30352) );
  OA22X1 U6698 ( .IN1(n4151), .IN2(n4152), .IN3(n1497), .IN4(n5626), .Q(n4149)
         );
  OA21X1 U6699 ( .IN1(n5460), .IN2(n4151), .IN3(n6408), .Q(n4150) );
  NAND2X0 U6700 ( .IN1(n5460), .IN2(n5780), .QN(n4152) );
  OAI22X1 U6701 ( .IN1(n4364), .IN2(n6145), .IN3(n4365), .IN4(n5781), .QN(
        g29260) );
  OA22X1 U6702 ( .IN1(n1589), .IN2(n4366), .IN3(n4363), .IN4(n5861), .Q(n4364)
         );
  OA21X1 U6703 ( .IN1(n1589), .IN2(n5423), .IN3(n6367), .Q(n4365) );
  NAND2X0 U6704 ( .IN1(n5423), .IN2(n5781), .QN(n4366) );
  OAI22X1 U6705 ( .IN1(n4077), .IN2(n6145), .IN3(n4078), .IN4(n5782), .QN(
        g30382) );
  OA22X1 U6706 ( .IN1(n4079), .IN2(n4080), .IN3(n1640), .IN4(n5625), .Q(n4077)
         );
  OA21X1 U6707 ( .IN1(n5461), .IN2(n4079), .IN3(n6405), .Q(n4078) );
  NAND2X0 U6708 ( .IN1(n5461), .IN2(n5782), .QN(n4080) );
  OAI22X1 U6709 ( .IN1(n6303), .IN2(n5769), .IN3(n2671), .IN4(n6141), .QN(
        g34264) );
  OA22X1 U6710 ( .IN1(n5613), .IN2(n2672), .IN3(n2673), .IN4(n1384), .Q(n2671)
         );
  INVX0 U6711 ( .IN(n2672), .QN(n1384) );
  NAND2X0 U6712 ( .IN1(n2675), .IN2(n2676), .QN(n2672) );
  OAI22X1 U6713 ( .IN1(n6300), .IN2(n5770), .IN3(n2650), .IN4(n6141), .QN(
        g34269) );
  OA22X1 U6714 ( .IN1(n5614), .IN2(n2651), .IN3(n2652), .IN4(n1389), .Q(n2650)
         );
  INVX0 U6715 ( .IN(n2651), .QN(n1389) );
  NAND2X0 U6716 ( .IN1(n2654), .IN2(n2655), .QN(n2651) );
  OAI22X1 U6717 ( .IN1(n6322), .IN2(n5577), .IN3(n5052), .IN4(n6141), .QN(
        g25636) );
  OA22X1 U6718 ( .IN1(n5381), .IN2(n5053), .IN3(n1549), .IN4(n5796), .Q(n5052)
         );
  INVX0 U6719 ( .IN(n5053), .QN(n1549) );
  NAND2X0 U6720 ( .IN1(n6024), .IN2(n2035), .QN(n5053) );
  OAI22X1 U6721 ( .IN1(n6318), .IN2(n5813), .IN3(n2926), .IN4(n6140), .QN(
        g33981) );
  OA22X1 U6722 ( .IN1(n2910), .IN2(n2927), .IN3(n1361), .IN4(n5793), .Q(n2926)
         );
  INVX0 U6723 ( .IN(n2927), .QN(n1361) );
  NAND2X0 U6724 ( .IN1(n2923), .IN2(n5534), .QN(n2927) );
  OAI22X1 U6725 ( .IN1(n6310), .IN2(n5815), .IN3(n2856), .IN4(n6142), .QN(
        g34002) );
  OA22X1 U6726 ( .IN1(n2839), .IN2(n2857), .IN3(n1322), .IN4(n5794), .Q(n2856)
         );
  INVX0 U6727 ( .IN(n2857), .QN(n1322) );
  NAND2X0 U6728 ( .IN1(n2853), .IN2(n5537), .QN(n2857) );
  OAI22X1 U6729 ( .IN1(n6314), .IN2(n5795), .IN3(n2941), .IN4(n6143), .QN(
        g33977) );
  OA22X1 U6730 ( .IN1(n2933), .IN2(n2942), .IN3(n1355), .IN4(n5804), .Q(n2941)
         );
  INVX0 U6731 ( .IN(n2942), .QN(n1355) );
  NAND2X0 U6732 ( .IN1(n2943), .IN2(n5504), .QN(n2942) );
  OAI22X1 U6733 ( .IN1(n6310), .IN2(n5788), .IN3(n2871), .IN4(n6142), .QN(
        g33998) );
  OA22X1 U6734 ( .IN1(n2862), .IN2(n2872), .IN3(n1317), .IN4(n5803), .Q(n2871)
         );
  INVX0 U6735 ( .IN(n2872), .QN(n1317) );
  NAND2X0 U6736 ( .IN1(n2873), .IN2(n5514), .QN(n2872) );
  OAI22X1 U6737 ( .IN1(n6307), .IN2(n5816), .IN3(n2809), .IN4(n6142), .QN(
        g34016) );
  OA22X1 U6738 ( .IN1(n2792), .IN2(n2810), .IN3(n1338), .IN4(n5787), .Q(n2809)
         );
  INVX0 U6739 ( .IN(n2810), .QN(n1338) );
  NAND2X0 U6740 ( .IN1(n2806), .IN2(n5521), .QN(n2810) );
  OAI22X1 U6741 ( .IN1(n6311), .IN2(n5812), .IN3(n2879), .IN4(n6143), .QN(
        g33995) );
  OA22X1 U6742 ( .IN1(n2862), .IN2(n2880), .IN3(n1314), .IN4(n5788), .Q(n2879)
         );
  INVX0 U6743 ( .IN(n2880), .QN(n1314) );
  NAND2X0 U6744 ( .IN1(n2876), .IN2(n5538), .QN(n2880) );
  OAI22X1 U6745 ( .IN1(n6308), .IN2(n5789), .IN3(n2825), .IN4(n6142), .QN(
        g34012) );
  OA22X1 U6746 ( .IN1(n2816), .IN2(n2826), .IN3(n1333), .IN4(n5798), .Q(n2825)
         );
  INVX0 U6747 ( .IN(n2826), .QN(n1333) );
  NAND2X0 U6748 ( .IN1(n2827), .IN2(n5523), .QN(n2826) );
  OAI22X1 U6749 ( .IN1(n6312), .IN2(n5818), .IN3(n2902), .IN4(n6142), .QN(
        g33988) );
  OA22X1 U6750 ( .IN1(n2886), .IN2(n2903), .IN3(n1370), .IN4(n5790), .Q(n2902)
         );
  INVX0 U6751 ( .IN(n2903), .QN(n1370) );
  NAND2X0 U6752 ( .IN1(n2899), .IN2(n5535), .QN(n2903) );
  OAI22X1 U6753 ( .IN1(n6309), .IN2(n5814), .IN3(n2833), .IN4(n6142), .QN(
        g34009) );
  OA22X1 U6754 ( .IN1(n2816), .IN2(n2834), .IN3(n1330), .IN4(n5789), .Q(n2833)
         );
  INVX0 U6755 ( .IN(n2834), .QN(n1330) );
  NAND2X0 U6756 ( .IN1(n2830), .IN2(n5522), .QN(n2834) );
  OAI22X1 U6757 ( .IN1(n6312), .IN2(n5790), .IN3(n2894), .IN4(n6143), .QN(
        g33991) );
  OA22X1 U6758 ( .IN1(n2886), .IN2(n2895), .IN3(n1373), .IN4(n5801), .Q(n2894)
         );
  INVX0 U6759 ( .IN(n2895), .QN(n1373) );
  NAND2X0 U6760 ( .IN1(n2896), .IN2(n5505), .QN(n2895) );
  OAI22X1 U6761 ( .IN1(n6318), .IN2(n5791), .IN3(n2967), .IN4(n6144), .QN(
        g33969) );
  OA22X1 U6762 ( .IN1(n2956), .IN2(n2968), .IN3(n1346), .IN4(n5587), .Q(n2967)
         );
  INVX0 U6763 ( .IN(n2968), .QN(n1346) );
  NAND2X0 U6764 ( .IN1(n2969), .IN2(n5362), .QN(n2968) );
  OAI22X1 U6765 ( .IN1(n6300), .IN2(n5811), .IN3(n2973), .IN4(n6141), .QN(
        g33967) );
  OA22X1 U6766 ( .IN1(n2956), .IN2(n2974), .IN3(n1345), .IN4(n5792), .Q(n2973)
         );
  INVX0 U6767 ( .IN(n2974), .QN(n1345) );
  NAND2X0 U6768 ( .IN1(n2969), .IN2(n5598), .QN(n2974) );
  OAI22X1 U6769 ( .IN1(n6313), .IN2(n5793), .IN3(n2918), .IN4(n6143), .QN(
        g33984) );
  OA22X1 U6770 ( .IN1(n2910), .IN2(n2919), .IN3(n1364), .IN4(n5799), .Q(n2918)
         );
  INVX0 U6771 ( .IN(n2919), .QN(n1364) );
  NAND2X0 U6772 ( .IN1(n2920), .IN2(n5503), .QN(n2919) );
  OAI22X1 U6773 ( .IN1(n6309), .IN2(n5794), .IN3(n2848), .IN4(n6143), .QN(
        g34005) );
  OA22X1 U6774 ( .IN1(n2839), .IN2(n2849), .IN3(n1325), .IN4(n5802), .Q(n2848)
         );
  INVX0 U6775 ( .IN(n2849), .QN(n1325) );
  NAND2X0 U6776 ( .IN1(n2850), .IN2(n5513), .QN(n2849) );
  OAI22X1 U6777 ( .IN1(n6315), .IN2(n5817), .IN3(n2949), .IN4(n6143), .QN(
        g33974) );
  OA22X1 U6778 ( .IN1(n2933), .IN2(n2950), .IN3(n1352), .IN4(n5795), .Q(n2949)
         );
  INVX0 U6779 ( .IN(n2950), .QN(n1352) );
  NAND2X0 U6780 ( .IN1(n2946), .IN2(n5536), .QN(n2950) );
  OAI22X1 U6781 ( .IN1(n6308), .IN2(n5798), .IN3(n2828), .IN4(n6142), .QN(
        g34011) );
  OA22X1 U6782 ( .IN1(n2816), .IN2(n2829), .IN3(n1331), .IN4(n5685), .Q(n2828)
         );
  INVX0 U6783 ( .IN(n2829), .QN(n1331) );
  NAND2X0 U6784 ( .IN1(n2830), .IN2(n5357), .QN(n2829) );
  OAI22X1 U6785 ( .IN1(n6313), .IN2(n5799), .IN3(n2921), .IN4(n6143), .QN(
        g33983) );
  OA22X1 U6786 ( .IN1(n2910), .IN2(n2922), .IN3(n1362), .IN4(n5686), .Q(n2921)
         );
  INVX0 U6787 ( .IN(n2922), .QN(n1362) );
  NAND2X0 U6788 ( .IN1(n2923), .IN2(n5354), .QN(n2922) );
  OAI22X1 U6789 ( .IN1(n6307), .IN2(n5800), .IN3(n2804), .IN4(n6141), .QN(
        g34018) );
  OA22X1 U6790 ( .IN1(n2792), .IN2(n2805), .IN3(n1339), .IN4(n5684), .Q(n2804)
         );
  INVX0 U6791 ( .IN(n2805), .QN(n1339) );
  NAND2X0 U6792 ( .IN1(n2806), .IN2(n5351), .QN(n2805) );
  OAI22X1 U6793 ( .IN1(n6305), .IN2(n5801), .IN3(n2897), .IN4(n6143), .QN(
        g33990) );
  OA22X1 U6794 ( .IN1(n2886), .IN2(n2898), .IN3(n1371), .IN4(n5683), .Q(n2897)
         );
  INVX0 U6795 ( .IN(n2898), .QN(n1371) );
  NAND2X0 U6796 ( .IN1(n2899), .IN2(n5355), .QN(n2898) );
  OAI22X1 U6797 ( .IN1(n6309), .IN2(n5802), .IN3(n2851), .IN4(n6143), .QN(
        g34004) );
  OA22X1 U6798 ( .IN1(n2839), .IN2(n2852), .IN3(n1323), .IN4(n5687), .Q(n2851)
         );
  INVX0 U6799 ( .IN(n2852), .QN(n1323) );
  NAND2X0 U6800 ( .IN1(n2853), .IN2(n5353), .QN(n2852) );
  OAI22X1 U6801 ( .IN1(n6311), .IN2(n5803), .IN3(n2874), .IN4(n6143), .QN(
        g33997) );
  OA22X1 U6802 ( .IN1(n2862), .IN2(n2875), .IN3(n1315), .IN4(n5688), .Q(n2874)
         );
  INVX0 U6803 ( .IN(n2875), .QN(n1315) );
  NAND2X0 U6804 ( .IN1(n2876), .IN2(n5356), .QN(n2875) );
  OAI22X1 U6805 ( .IN1(n6314), .IN2(n5804), .IN3(n2944), .IN4(n6143), .QN(
        g33976) );
  OA22X1 U6806 ( .IN1(n2933), .IN2(n2945), .IN3(n1353), .IN4(n5797), .Q(n2944)
         );
  INVX0 U6807 ( .IN(n2945), .QN(n1353) );
  NAND2X0 U6808 ( .IN1(n2946), .IN2(n5352), .QN(n2945) );
  NAND2X0 U6809 ( .IN1(n6232), .IN2(n5714), .QN(n4865) );
  NAND2X0 U6810 ( .IN1(n3005), .IN2(n5359), .QN(n3002) );
  INVX0 U6811 ( .IN(n4853), .QN(n1426) );
  INVX0 U6812 ( .IN(n4852), .QN(n1427) );
  AO21X1 U6813 ( .IN1(n4062), .IN2(n4444), .IN3(n4051), .Q(n3610) );
  NAND2X0 U6814 ( .IN1(n4388), .IN2(n5403), .QN(n4444) );
  AO21X1 U6815 ( .IN1(n4062), .IN2(n4399), .IN3(n4051), .Q(n3535) );
  NAND2X0 U6816 ( .IN1(n4388), .IN2(n5404), .QN(n4399) );
  INVX0 U6817 ( .IN(n5027), .QN(n1436) );
  INVX0 U6818 ( .IN(g34025), .QN(n1297) );
  INVX0 U6819 ( .IN(n3338), .QN(n1793) );
  INVX0 U6820 ( .IN(n2760), .QN(n1300) );
  INVX0 U6821 ( .IN(n3146), .QN(n1483) );
  INVX0 U6822 ( .IN(n4139), .QN(n1852) );
  INVX0 U6823 ( .IN(n4091), .QN(n1742) );
  INVX0 U6824 ( .IN(n3206), .QN(n1479) );
  INVX0 U6825 ( .IN(n3226), .QN(n1477) );
  INVX0 U6826 ( .IN(n3186), .QN(n1481) );
  INVX0 U6827 ( .IN(n3748), .QN(n1516) );
  INVX0 U6828 ( .IN(n4147), .QN(n1853) );
  INVX0 U6829 ( .IN(n4099), .QN(n1743) );
  NAND4X0 U6830 ( .IN1(n4800), .IN2(n4801), .IN3(n4802), .IN4(n5466), .QN(
        n3258) );
  NAND4X0 U6831 ( .IN1(n4807), .IN2(n4808), .IN3(n4809), .IN4(n5467), .QN(
        n3266) );
  NOR2X0 U6832 ( .IN1(n4340), .IN2(n3069), .QN(n4333) );
  NOR2X0 U6833 ( .IN1(n4234), .IN2(n3027), .QN(n4227) );
  NOR2X0 U6834 ( .IN1(n4279), .IN2(n1560), .QN(n4272) );
  NOR2X0 U6835 ( .IN1(n4264), .IN2(n1562), .QN(n4257) );
  NOR2X0 U6836 ( .IN1(n4219), .IN2(n1705), .QN(n4212) );
  NOR2X0 U6837 ( .IN1(n4370), .IN2(n1590), .QN(n4363) );
  NOR2X0 U6838 ( .IN1(n4355), .IN2(n1650), .QN(n4348) );
  NOR2X0 U6839 ( .IN1(n4249), .IN2(n1564), .QN(n4242) );
  NOR2X0 U6840 ( .IN1(n5160), .IN2(n5515), .QN(n5158) );
  NOR2X0 U6841 ( .IN1(n5155), .IN2(n5529), .QN(n5153) );
  NOR2X0 U6842 ( .IN1(n5140), .IN2(n5531), .QN(n5138) );
  NOR2X0 U6843 ( .IN1(n5150), .IN2(n5528), .QN(n5148) );
  NOR2X0 U6844 ( .IN1(n5182), .IN2(n5530), .QN(n5180) );
  NOR2X0 U6845 ( .IN1(n5145), .IN2(n5533), .QN(n5143) );
  NOR2X0 U6846 ( .IN1(n5192), .IN2(n5527), .QN(n5190) );
  NOR2X0 U6847 ( .IN1(n5187), .IN2(n5532), .QN(n5185) );
  NAND2X0 U6848 ( .IN1(n5386), .IN2(n5563), .QN(n3773) );
  NAND2X0 U6849 ( .IN1(n5383), .IN2(n5569), .QN(n3983) );
  NAND2X0 U6850 ( .IN1(n5385), .IN2(n5568), .QN(n3807) );
  NAND2X0 U6851 ( .IN1(n5384), .IN2(n5567), .QN(n3907) );
  NAND2X0 U6852 ( .IN1(n5389), .IN2(n5566), .QN(n3874) );
  NAND2X0 U6853 ( .IN1(n5387), .IN2(n5564), .QN(n3950) );
  NAND2X0 U6854 ( .IN1(n5388), .IN2(n5565), .QN(n3841) );
  NAND2X0 U6855 ( .IN1(n5603), .IN2(n5390), .QN(n4014) );
  NAND2X0 U6856 ( .IN1(n5067), .IN2(n4176), .QN(n5063) );
  NAND2X0 U6857 ( .IN1(n5319), .IN2(n5616), .QN(n4176) );
  NAND2X0 U6858 ( .IN1(n5320), .IN2(n5622), .QN(n4194) );
  NAND2X0 U6859 ( .IN1(n3706), .IN2(n5578), .QN(n3698) );
  NAND2X0 U6860 ( .IN1(n2751), .IN2(n2669), .QN(n2755) );
  NAND2X0 U6861 ( .IN1(n2766), .IN2(n2689), .QN(n2770) );
  NAND4X0 U6862 ( .IN1(n5628), .IN2(n5413), .IN3(n5315), .IN4(n5280), .QN(
        n2442) );
  NAND2X0 U6863 ( .IN1(n5067), .IN2(n5322), .QN(n4801) );
  NAND2X0 U6864 ( .IN1(n2582), .IN2(n5382), .QN(n2579) );
  NAND2X0 U6865 ( .IN1(n5480), .IN2(n5340), .QN(n3286) );
  NAND2X0 U6866 ( .IN1(n5400), .IN2(n5604), .QN(n4687) );
  NAND2X0 U6867 ( .IN1(n5588), .IN2(n5393), .QN(n4658) );
  NAND2X0 U6868 ( .IN1(n5589), .IN2(n5394), .QN(n4612) );
  NAND2X0 U6869 ( .IN1(n5593), .IN2(n5397), .QN(n4635) );
  NAND2X0 U6870 ( .IN1(n5594), .IN2(n5395), .QN(n4677) );
  NAND2X0 U6871 ( .IN1(n5590), .IN2(n5398), .QN(n4566) );
  NAND2X0 U6872 ( .IN1(n5591), .IN2(n5399), .QN(n4682) );
  NAND2X0 U6873 ( .IN1(n5592), .IN2(n5396), .QN(n4589) );
  NAND2X0 U6874 ( .IN1(n2604), .IN2(n2582), .QN(n2596) );
  NAND2X0 U6875 ( .IN1(n3115), .IN2(n1474), .QN(n3242) );
  NAND2X0 U6876 ( .IN1(n3115), .IN2(n1482), .QN(n3162) );
  NAND2X0 U6877 ( .IN1(n3115), .IN2(n1481), .QN(n3183) );
  NAND2X0 U6878 ( .IN1(n3115), .IN2(n1477), .QN(n3223) );
  NAND2X0 U6879 ( .IN1(n3115), .IN2(n1483), .QN(n3143) );
  NAND2X0 U6880 ( .IN1(n3115), .IN2(n1479), .QN(n3203) );
  NAND2X0 U6881 ( .IN1(n2675), .IN2(n2688), .QN(n2686) );
  NAND2X0 U6882 ( .IN1(n2654), .IN2(n2667), .QN(n2665) );
  NAND2X0 U6883 ( .IN1(n2654), .IN2(n2659), .QN(n2657) );
  NAND2X0 U6884 ( .IN1(n2675), .IN2(n2680), .QN(n2678) );
  NAND2X0 U6885 ( .IN1(n3833), .IN2(n1843), .QN(n3429) );
  NAND2X0 U6886 ( .IN1(n3833), .IN2(n1842), .QN(n3409) );
  NAND2X0 U6887 ( .IN1(n2675), .IN2(n2684), .QN(n2682) );
  NAND2X0 U6888 ( .IN1(n2654), .IN2(n2663), .QN(n2661) );
  NAND2X0 U6889 ( .IN1(n3833), .IN2(n1845), .QN(n3419) );
  NAND2X0 U6890 ( .IN1(n3833), .IN2(n1844), .QN(n3439) );
  NAND2X0 U6891 ( .IN1(n2669), .IN2(n2670), .QN(n2560) );
  NAND2X0 U6892 ( .IN1(n2689), .IN2(n2690), .QN(n2570) );
  NAND3X0 U6893 ( .IN1(n3282), .IN2(n2515), .IN3(n2714), .QN(g33659) );
  NOR2X0 U6894 ( .IN1(n4052), .IN2(n5301), .QN(n4064) );
  AND3X1 U6895 ( .IN1(n3023), .IN2(n1484), .IN3(n3088), .Q(n3086) );
  NAND2X0 U6896 ( .IN1(n1987), .IN2(n5321), .QN(n4808) );
  NOR4X0 U6897 ( .IN1(n3719), .IN2(n3720), .IN3(n3721), .IN4(n3722), .QN(n3712) );
  AND3X1 U6898 ( .IN1(n3023), .IN2(n1487), .IN3(g28753), .Q(n3052) );
  NAND3X0 U6899 ( .IN1(n3653), .IN2(n5600), .IN3(n4062), .QN(n4050) );
  NAND3X0 U6900 ( .IN1(n5518), .IN2(n5361), .IN3(n1558), .QN(n2684) );
  NAND3X0 U6901 ( .IN1(n5517), .IN2(n5360), .IN3(n1704), .QN(n2663) );
  AND3X1 U6902 ( .IN1(n3033), .IN2(n1486), .IN3(n3079), .Q(n3075) );
  AND3X1 U6903 ( .IN1(n3023), .IN2(n1486), .IN3(n3018), .Q(n3014) );
  AND3X1 U6904 ( .IN1(n3033), .IN2(n1487), .IN3(n3038), .Q(n3034) );
  AND3X1 U6905 ( .IN1(n3023), .IN2(n1488), .IN3(n3047), .Q(n3043) );
  AND3X1 U6906 ( .IN1(n5607), .IN2(n5950), .IN3(n4670), .Q(n3720) );
  NAND2X0 U6907 ( .IN1(g27831), .IN2(n3240), .QN(n3243) );
  AND3X1 U6908 ( .IN1(n5711), .IN2(n5416), .IN3(n4724), .Q(n4726) );
  AND3X1 U6909 ( .IN1(n5543), .IN2(n5350), .IN3(n1844), .Q(n4725) );
  AO21X1 U6910 ( .IN1(n5327), .IN2(n4828), .IN3(n4829), .Q(n4542) );
  ISOLANDX1 U6911 ( .D(n3115), .ISO(n2726), .Q(n3111) );
  ISOLANDX1 U6912 ( .D(n3115), .ISO(n2727), .Q(n3131) );
  INVX0 U6913 ( .IN(g28753), .QN(n1560) );
  NOR2X0 U6914 ( .IN1(n2631), .IN2(n2632), .QN(n2612) );
  NOR2X0 U6915 ( .IN1(n2637), .IN2(n2631), .QN(n2622) );
  NOR2X0 U6916 ( .IN1(n2048), .IN2(n2631), .QN(n2626) );
  ISOLANDX1 U6917 ( .D(n3933), .ISO(n5350), .Q(n3799) );
  INVX0 U6918 ( .IN(n3287), .QN(g32975) );
  INVX0 U6919 ( .IN(g27831), .QN(n1599) );
  NOR2X0 U6920 ( .IN1(n3729), .IN2(n5340), .QN(n3472) );
  NOR2X0 U6921 ( .IN1(n5612), .IN2(n4723), .QN(n4729) );
  INVX0 U6922 ( .IN(n2724), .QN(g31862) );
  NOR2X0 U6923 ( .IN1(n5543), .IN2(n4328), .QN(n3942) );
  INVX0 U6924 ( .IN(n2739), .QN(g31860) );
  NOR2X0 U6925 ( .IN1(n2604), .IN2(n5539), .QN(n2601) );
  ISOLANDX1 U6926 ( .D(n3664), .ISO(n5674), .Q(n3662) );
  ISOLANDX1 U6927 ( .D(n3673), .ISO(n5673), .Q(n3671) );
  NOR2X0 U6928 ( .IN1(n2609), .IN2(n5348), .QN(n2607) );
  ISOLANDX1 U6929 ( .D(n3505), .ISO(n3506), .Q(n2790) );
  OR2X1 U6930 ( .IN1(n2693), .IN2(n5298), .Q(n2609) );
  ISOLANDX1 U6931 ( .D(n4490), .ISO(n5554), .Q(n4178) );
  ISOLANDX1 U6932 ( .D(n4514), .ISO(n5555), .Q(n4196) );
  ISOLANDX1 U6933 ( .D(n4178), .ISO(n5558), .Q(n3736) );
  ISOLANDX1 U6934 ( .D(n4196), .ISO(n5559), .Q(n3741) );
  ISOLANDX1 U6935 ( .D(n3736), .ISO(n5553), .Q(n3664) );
  ISOLANDX1 U6936 ( .D(n3741), .ISO(n5560), .Q(n3673) );
  ISOLANDX1 U6937 ( .D(n2601), .ISO(n5303), .Q(n2598) );
  ISOLANDX1 U6938 ( .D(n4804), .ISO(n5556), .Q(n4490) );
  ISOLANDX1 U6939 ( .D(n4811), .ISO(n5557), .Q(n4514) );
  ISOLANDX1 U6940 ( .D(n4814), .ISO(n5422), .Q(n4519) );
  ISOLANDX1 U6941 ( .D(n2607), .ISO(n5323), .Q(n2594) );
  NAND3X0 U6942 ( .IN1(n5304), .IN2(n5622), .IN3(n5392), .QN(n5084) );
  NAND3X0 U6943 ( .IN1(n5401), .IN2(n5302), .IN3(n5616), .QN(n5060) );
  ISOLANDX1 U6944 ( .D(n3084), .ISO(n5348), .Q(n3033) );
  NAND2X0 U6945 ( .IN1(n4295), .IN2(n3013), .QN(n4692) );
  NAND2X0 U6946 ( .IN1(n4317), .IN2(n3012), .QN(n4698) );
  NOR2X0 U6947 ( .IN1(n2076), .IN2(n5709), .QN(n4953) );
  INVX0 U6948 ( .IN(n3004), .QN(g31863) );
  NAND2X0 U6949 ( .IN1(n6022), .IN2(n3510), .QN(n3512) );
  ISOLANDX1 U6950 ( .D(n2598), .ISO(n5365), .Q(n2590) );
  OR3X1 U6951 ( .IN1(n5067), .IN2(n5066), .IN3(n5322), .Q(n4802) );
  OR3X1 U6952 ( .IN1(n1987), .IN2(n5090), .IN3(n5321), .Q(n4809) );
  AND2X1 U6953 ( .IN1(n4724), .IN2(n4725), .Q(n4722) );
  ISOLANDX1 U6954 ( .D(n3122), .ISO(n2727), .Q(n3125) );
  ISOLANDX1 U6955 ( .D(n3102), .ISO(n2726), .Q(n3105) );
  ISOLANDX1 U6956 ( .D(n3141), .ISO(n3146), .Q(n3145) );
  ISOLANDX1 U6957 ( .D(n3160), .ISO(n3165), .Q(n3164) );
  AO21X1 U6958 ( .IN1(n2417), .IN2(n5653), .IN3(n5298), .Q(n2409) );
  NAND2X0 U6959 ( .IN1(n3621), .IN2(n6022), .QN(n3623) );
  OA22X1 U6960 ( .IN1(n3291), .IN2(n3298), .IN3(n3293), .IN4(n3299), .Q(n3297)
         );
  OA22X1 U6961 ( .IN1(n3291), .IN2(n3292), .IN3(n3293), .IN4(n3294), .Q(n3290)
         );
  OA21X1 U6962 ( .IN1(n1381), .IN2(n5771), .IN3(n2674), .Q(n2687) );
  OA21X1 U6963 ( .IN1(n1381), .IN2(n5769), .IN3(n2674), .Q(n2673) );
  OA21X1 U6964 ( .IN1(n1386), .IN2(n5770), .IN3(n2653), .Q(n2652) );
  OA21X1 U6965 ( .IN1(n1386), .IN2(n5772), .IN3(n2653), .Q(n2658) );
  OA21X1 U6966 ( .IN1(n1381), .IN2(n5773), .IN3(n2674), .Q(n2683) );
  OA21X1 U6967 ( .IN1(n1386), .IN2(n5774), .IN3(n2653), .Q(n2666) );
  OA21X1 U6968 ( .IN1(n1381), .IN2(n5775), .IN3(n2674), .Q(n2679) );
  OA21X1 U6969 ( .IN1(n1386), .IN2(n5776), .IN3(n2653), .Q(n2662) );
  NAND2X0 U6970 ( .IN1(n3547), .IN2(n6022), .QN(n3549) );
  NAND2X0 U6971 ( .IN1(n3585), .IN2(n6022), .QN(n3587) );
  NAND2X0 U6972 ( .IN1(n3603), .IN2(n6022), .QN(n3605) );
  NAND2X0 U6973 ( .IN1(n3529), .IN2(n6022), .QN(n3531) );
  NAND2X0 U6974 ( .IN1(n3566), .IN2(n6022), .QN(n3568) );
  NAND2X0 U6975 ( .IN1(n3639), .IN2(n6022), .QN(n3641) );
  NOR2X0 U6976 ( .IN1(n3206), .IN2(n1602), .QN(n3205) );
  NOR2X0 U6977 ( .IN1(n3226), .IN2(n1601), .QN(n3225) );
  NOR2X0 U6978 ( .IN1(n3186), .IN2(n1600), .QN(n3185) );
  NOR3X0 U6979 ( .IN1(n3235), .IN2(n4919), .IN3(n5304), .QN(n4184) );
  NOR3X0 U6980 ( .IN1(n3155), .IN2(n4894), .IN3(n5302), .QN(n4166) );
  NAND2X0 U6981 ( .IN1(n3688), .IN2(n5611), .QN(n3711) );
  INVX0 U6982 ( .IN(n4532), .QN(n1538) );
  OR2X1 U6983 ( .IN1(n2784), .IN2(n1490), .Q(n2782) );
  INVX0 U6984 ( .IN(n3088), .QN(n1590) );
  INVX0 U6985 ( .IN(n3079), .QN(n1650) );
  INVX0 U6986 ( .IN(n3018), .QN(n1705) );
  INVX0 U6987 ( .IN(n3047), .QN(n1562) );
  INVX0 U6988 ( .IN(n3038), .QN(n1564) );
  NAND2X0 U6989 ( .IN1(n3201), .IN2(n3202), .QN(n3204) );
  NAND2X0 U6990 ( .IN1(n3221), .IN2(n3222), .QN(n3224) );
  INVX0 U6991 ( .IN(n5226), .QN(n1740) );
  INVX0 U6992 ( .IN(n5204), .QN(n1570) );
  NAND2X0 U6993 ( .IN1(n3181), .IN2(n3182), .QN(n3184) );
  INVX0 U6994 ( .IN(n4052), .QN(n2138) );
  INVX0 U6995 ( .IN(n3027), .QN(n1565) );
  INVX0 U6996 ( .IN(n3069), .QN(n1611) );
  INVX0 U6997 ( .IN(n2582), .QN(n1299) );
  INVX0 U6998 ( .IN(n4504), .QN(n1693) );
  INVX0 U6999 ( .IN(n4480), .QN(n1776) );
  INVX0 U7000 ( .IN(n4051), .QN(n2140) );
  INVX0 U7001 ( .IN(n3296), .QN(n1546) );
  INVX0 U7002 ( .IN(n3910), .QN(n1581) );
  INVX0 U7003 ( .IN(n3776), .QN(n2224) );
  INVX0 U7004 ( .IN(n3877), .QN(n1968) );
  INVX0 U7005 ( .IN(n3810), .QN(n1514) );
  INVX0 U7006 ( .IN(n4017), .QN(n1730) );
  INVX0 U7007 ( .IN(n3953), .QN(n1908) );
  INVX0 U7008 ( .IN(n3986), .QN(n1680) );
  INVX0 U7009 ( .IN(n3844), .QN(n1821) );
  INVX0 U7010 ( .IN(n5094), .QN(n1987) );
  INVX0 U7011 ( .IN(n3288), .QN(n1843) );
  INVX0 U7012 ( .IN(n3201), .QN(n1602) );
  INVX0 U7013 ( .IN(n3289), .QN(n1755) );
  INVX0 U7014 ( .IN(n3295), .QN(n2223) );
  INVX0 U7015 ( .IN(n3221), .QN(n1601) );
  INVX0 U7016 ( .IN(n3298), .QN(n1907) );
  INVX0 U7017 ( .IN(n3292), .QN(n1513) );
  INVX0 U7018 ( .IN(n3294), .QN(n1820) );
  INVX0 U7019 ( .IN(n3299), .QN(n1679) );
  INVX0 U7020 ( .IN(n3181), .QN(n1600) );
  NAND2X0 U7021 ( .IN1(n3122), .IN2(n3123), .QN(n3124) );
  NAND2X0 U7022 ( .IN1(n5518), .IN2(n5361), .QN(n4325) );
  NAND2X0 U7023 ( .IN1(n5517), .IN2(n5360), .QN(n4303) );
  INVX0 U7024 ( .IN(n2750), .QN(n2136) );
  INVX0 U7025 ( .IN(n2765), .QN(n2103) );
  INVX0 U7026 ( .IN(n3634), .QN(n1952) );
  INVX0 U7027 ( .IN(n3235), .QN(n1696) );
  NAND2X0 U7028 ( .IN1(n3141), .IN2(n3142), .QN(n3144) );
  NAND2X0 U7029 ( .IN1(n3160), .IN2(n3161), .QN(n3163) );
  NAND2X0 U7030 ( .IN1(n3102), .IN2(n3103), .QN(n3104) );
  INVX0 U7031 ( .IN(n3291), .QN(n1842) );
  INVX0 U7032 ( .IN(n3293), .QN(n1845) );
  INVX0 U7033 ( .IN(n3155), .QN(n2034) );
  INVX0 U7034 ( .IN(n2741), .QN(n1880) );
  INVX0 U7035 ( .IN(n3659), .QN(n1572) );
  INVX0 U7036 ( .IN(n3668), .QN(n1582) );
  INVX0 U7037 ( .IN(n3706), .QN(n1809) );
  INVX0 U7038 ( .IN(n3705), .QN(n1823) );
  INVX0 U7039 ( .IN(n3090), .QN(n1881) );
  INVX0 U7040 ( .IN(n2675), .QN(n1381) );
  INVX0 U7041 ( .IN(n2654), .QN(n1386) );
  INVX0 U7042 ( .IN(n3056), .QN(n1893) );
  INVX0 U7043 ( .IN(n3019), .QN(n2122) );
  INVX0 U7044 ( .IN(n3039), .QN(n1869) );
  INVX0 U7045 ( .IN(n3080), .QN(n1941) );
  INVX0 U7046 ( .IN(n3029), .QN(n1624) );
  INVX0 U7047 ( .IN(n3048), .QN(n2304) );
  INVX0 U7048 ( .IN(n3071), .QN(n1749) );
  INVX0 U7049 ( .IN(n2736), .QN(n2123) );
  INVX0 U7050 ( .IN(n2743), .QN(n1940) );
  INVX0 U7051 ( .IN(n2734), .QN(n2307) );
  INVX0 U7052 ( .IN(n2742), .QN(n1625) );
  INVX0 U7053 ( .IN(n2745), .QN(n1870) );
  INVX0 U7054 ( .IN(n2746), .QN(n1747) );
  INVX0 U7055 ( .IN(n2752), .QN(n2135) );
  INVX0 U7056 ( .IN(n2767), .QN(n2101) );
  INVX0 U7057 ( .IN(n3215), .QN(n1694) );
  NAND2X0 U7058 ( .IN1(n4317), .IN2(n4318), .QN(n4311) );
  XNOR2X1 U7059 ( .IN1(n4319), .IN2(g34657), .Q(n4318) );
  OA221X1 U7060 ( .IN1(n5344), .IN2(n2765), .IN3(n5296), .IN4(n2767), .IN5(
        n4324), .Q(n4319) );
  OA22X1 U7061 ( .IN1(n5345), .IN2(n4325), .IN3(n5312), .IN4(n4326), .Q(n4324)
         );
  NAND2X0 U7062 ( .IN1(n4295), .IN2(n4296), .QN(n4289) );
  XNOR2X1 U7063 ( .IN1(n4297), .IN2(g34649), .Q(n4296) );
  OA221X1 U7064 ( .IN1(n5295), .IN2(n2750), .IN3(n5346), .IN4(n2752), .IN5(
        n4302), .Q(n4297) );
  OA22X1 U7065 ( .IN1(n5297), .IN2(n4303), .IN3(n5408), .IN4(n4304), .Q(n4302)
         );
  INVX0 U7066 ( .IN(n3135), .QN(n2035) );
  INVX0 U7067 ( .IN(n2754), .QN(n1608) );
  INVX0 U7068 ( .IN(n2769), .QN(n1727) );
  INVX0 U7069 ( .IN(n3599), .QN(n2228) );
  INVX0 U7070 ( .IN(n3617), .QN(n1661) );
  INVX0 U7071 ( .IN(n3542), .QN(n2072) );
  INVX0 U7072 ( .IN(n3561), .QN(n1759) );
  INVX0 U7073 ( .IN(n3523), .QN(n1670) );
  INVX0 U7074 ( .IN(n3580), .QN(n2131) );
  INVX0 U7075 ( .IN(n3089), .QN(n1882) );
  INVX0 U7076 ( .IN(n2457), .QN(n2172) );
  INVX0 U7077 ( .IN(n3652), .QN(n2218) );
  INVX0 U7078 ( .IN(n3055), .QN(n1891) );
  INVX0 U7079 ( .IN(n3037), .QN(n1867) );
  INVX0 U7080 ( .IN(n3046), .QN(n2303) );
  INVX0 U7081 ( .IN(n3070), .QN(n1751) );
  INVX0 U7082 ( .IN(n3017), .QN(n2120) );
  INVX0 U7083 ( .IN(n3078), .QN(n1942) );
  INVX0 U7084 ( .IN(n3028), .QN(n1622) );
  INVX0 U7085 ( .IN(n3697), .QN(n1822) );
  INVX0 U7086 ( .IN(n4818), .QN(n2075) );
  INVX0 U7087 ( .IN(n2428), .QN(n1485) );
  INVX0 U7088 ( .IN(n3471), .QN(n1645) );
  INVX0 U7089 ( .IN(n4499), .QN(n1695) );
  INVX0 U7090 ( .IN(n4948), .QN(n2076) );
  INVX0 U7091 ( .IN(n2417), .QN(n1390) );
  INVX0 U7092 ( .IN(n2733), .QN(n1488) );
  INVX0 U7093 ( .IN(n2740), .QN(n1484) );
  INVX0 U7094 ( .IN(n2669), .QN(n1307) );
  INVX0 U7095 ( .IN(n2689), .QN(n1303) );
  INVX0 U7096 ( .IN(n4067), .QN(n1712) );
  INVX0 U7097 ( .IN(n4115), .QN(n1856) );
  INVX0 U7098 ( .IN(n4079), .QN(n1640) );
  INVX0 U7099 ( .IN(n4127), .QN(n1612) );
  INVX0 U7100 ( .IN(n4103), .QN(n1860) );
  INVX0 U7101 ( .IN(n4151), .QN(n1497) );
  INVX0 U7102 ( .IN(n3710), .QN(n1824) );
  INVX0 U7103 ( .IN(n4485), .QN(n1775) );
  INVX0 U7104 ( .IN(n4509), .QN(n1692) );
  INVX0 U7105 ( .IN(n4203), .QN(n1605) );
  INVX0 U7106 ( .IN(n3506), .QN(n2049) );
  INVX0 U7107 ( .IN(n3692), .QN(n1874) );
  INVX0 U7108 ( .IN(n4123), .QN(n1857) );
  INVX0 U7109 ( .IN(n4075), .QN(n1668) );
  INVX0 U7110 ( .IN(n4087), .QN(n1641) );
  INVX0 U7111 ( .IN(n4135), .QN(n1613) );
  INVX0 U7112 ( .IN(n4111), .QN(n1861) );
  INVX0 U7113 ( .IN(n4829), .QN(n1888) );
  INVX0 U7114 ( .IN(g24167), .QN(n1492) );
  INVX0 U7115 ( .IN(n2716), .QN(n1480) );
  INVX0 U7116 ( .IN(n2715), .QN(n1478) );
  INVX0 U7117 ( .IN(n2515), .QN(n1473) );
  INVX0 U7118 ( .IN(n2725), .QN(n1476) );
  NOR2X0 U7119 ( .IN1(n3770), .IN2(n5646), .QN(n3400) );
  NOR2X0 U7120 ( .IN1(n3904), .IN2(n5650), .QN(n3440) );
  NOR2X0 U7121 ( .IN1(n3804), .IN2(n5651), .QN(n3410) );
  NOR2X0 U7122 ( .IN1(n3947), .IN2(n5648), .QN(n3475) );
  NOR2X0 U7123 ( .IN1(n3838), .IN2(n5649), .QN(n3420) );
  NOR2X0 U7124 ( .IN1(n3871), .IN2(n5647), .QN(n3430) );
  NOR2X0 U7125 ( .IN1(n3980), .IN2(n5645), .QN(n3485) );
  NOR2X0 U7126 ( .IN1(n5768), .IN2(n5049), .QN(n5047) );
  NOR2X0 U7127 ( .IN1(n5767), .IN2(n5075), .QN(n5073) );
  INVX0 U7128 ( .IN(n4020), .QN(n1732) );
  INVX0 U7129 ( .IN(n3495), .QN(n1729) );
  INVX0 U7130 ( .IN(n3945), .QN(n1905) );
  INVX0 U7131 ( .IN(n3836), .QN(n1818) );
  INVX0 U7132 ( .IN(n3768), .QN(n2222) );
  INVX0 U7133 ( .IN(n3869), .QN(n1967) );
  INVX0 U7134 ( .IN(n3978), .QN(n1678) );
  INVX0 U7135 ( .IN(n3802), .QN(n1511) );
  INVX0 U7136 ( .IN(n3902), .QN(n1578) );
  INVX0 U7137 ( .IN(n3904), .QN(n1576) );
  INVX0 U7138 ( .IN(n3947), .QN(n1903) );
  INVX0 U7139 ( .IN(n3838), .QN(n1816) );
  INVX0 U7140 ( .IN(n3770), .QN(n2226) );
  INVX0 U7141 ( .IN(n3804), .QN(n1509) );
  INVX0 U7142 ( .IN(n3980), .QN(n1682) );
  INVX0 U7143 ( .IN(n3871), .QN(n1970) );
  INVX0 U7144 ( .IN(n4899), .QN(n1655) );
  INVX0 U7145 ( .IN(n4971), .QN(n1540) );
  INVX0 U7146 ( .IN(n4924), .QN(n1606) );
  NAND2X0 U7147 ( .IN1(n5463), .IN2(n5784), .QN(n4116) );
  NAND2X0 U7148 ( .IN1(n5464), .IN2(n5785), .QN(n4140) );
  NAND2X0 U7149 ( .IN1(n5424), .IN2(n5786), .QN(n4351) );
  NAND2X0 U7150 ( .IN1(n5462), .IN2(n5783), .QN(n4128) );
  NAND2X0 U7151 ( .IN1(n5425), .IN2(n5805), .QN(n4260) );
  NAND2X0 U7152 ( .IN1(n5426), .IN2(n5806), .QN(n4215) );
  NAND2X0 U7153 ( .IN1(n5427), .IN2(n5807), .QN(n4275) );
  NAND2X0 U7154 ( .IN1(n5428), .IN2(n5808), .QN(n4336) );
  NAND2X0 U7155 ( .IN1(n5429), .IN2(n5809), .QN(n4245) );
  NAND2X0 U7156 ( .IN1(n5430), .IN2(n5810), .QN(n4230) );
  INVX0 U7157 ( .IN(n5131), .QN(n1989) );
  INVX0 U7158 ( .IN(n4880), .QN(n1532) );
  AND3X1 U7159 ( .IN1(g562), .IN2(n4959), .IN3(n4960), .Q(n4826) );
  AO222X1 U7160 ( .IN1(n2649), .IN2(n5473), .IN3(n2705), .IN4(n2421), .IN5(
        g599), .IN6(n6094), .Q(g34251) );
  NOR2X0 U7161 ( .IN1(n2649), .IN2(n5473), .QN(n2705) );
  AO222X1 U7162 ( .IN1(n2423), .IN2(n5288), .IN3(n2426), .IN4(n2421), .IN5(
        g622), .IN6(n6096), .Q(g34849) );
  NOR2X0 U7163 ( .IN1(n2423), .IN2(n5288), .QN(n2426) );
  AO222X1 U7164 ( .IN1(n2509), .IN2(n5474), .IN3(n2555), .IN4(n2421), .IN5(
        g608), .IN6(n6097), .Q(g34599) );
  NOR2X0 U7165 ( .IN1(n2509), .IN2(n5474), .QN(n2555) );
  AO222X1 U7166 ( .IN1(n2487), .IN2(n5339), .IN3(n2508), .IN4(n2421), .IN5(
        g613), .IN6(n6094), .Q(g34724) );
  NOR2X0 U7167 ( .IN1(n2487), .IN2(n5339), .QN(n2508) );
  AO222X1 U7168 ( .IN1(n2427), .IN2(n5672), .IN3(n2486), .IN4(n2421), .IN5(
        g617), .IN6(n6095), .Q(g34790) );
  NOR2X0 U7169 ( .IN1(n2427), .IN2(n5672), .QN(n2486) );
  AO222X1 U7170 ( .IN1(n2556), .IN2(n5475), .IN3(n2648), .IN4(n2421), .IN5(
        g604), .IN6(n6092), .Q(g34438) );
  NOR2X0 U7171 ( .IN1(n2556), .IN2(n5475), .QN(n2648) );
  AO222X1 U7172 ( .IN1(n2420), .IN2(n2421), .IN3(n2422), .IN4(n5338), .IN5(
        g626), .IN6(n6096), .Q(g34880) );
  NOR2X0 U7173 ( .IN1(n2422), .IN2(n5338), .QN(n2420) );
  ISOLANDX1 U7174 ( .D(n2423), .ISO(n5288), .Q(n2422) );
  OR2X1 U7175 ( .IN1(g4405), .IN2(n5965), .Q(g26948) );
  AND3X1 U7176 ( .IN1(n4863), .IN2(n1648), .IN3(g4388), .Q(n5965) );
  AO221X1 U7177 ( .IN1(n2140), .IN2(n6152), .IN3(g2715), .IN4(n6087), .IN5(
        n5045), .Q(g25639) );
  AO22X1 U7178 ( .IN1(g559), .IN2(n6128), .IN3(n5114), .IN4(n2421), .Q(g25613)
         );
  OA21X1 U7179 ( .IN1(n5338), .IN2(n5288), .IN3(n5115), .Q(n5114) );
  XOR2X1 U7180 ( .IN1(g562), .IN2(n4960), .Q(n5115) );
  OR4X1 U7181 ( .IN1(g4411), .IN2(g7257), .IN3(g7243), .IN4(n5966), .Q(n4872)
         );
  OR2X1 U7182 ( .IN1(g4405), .IN2(g4375), .Q(n5966) );
  OA21X1 U7183 ( .IN1(n5485), .IN2(g9048), .IN3(g20763), .Q(n4960) );
  AO222X1 U7184 ( .IN1(n3684), .IN2(n5552), .IN3(n3744), .IN4(n2421), .IN5(
        g577), .IN6(n6102), .Q(g31866) );
  NOR2X0 U7185 ( .IN1(n3684), .IN2(n5552), .QN(n3744) );
  AO222X1 U7186 ( .IN1(n2706), .IN2(n5550), .IN3(n2981), .IN4(n2421), .IN5(
        g595), .IN6(n6100), .Q(g33964) );
  NOR2X0 U7187 ( .IN1(n2706), .IN2(n5550), .QN(n2981) );
  AO222X1 U7188 ( .IN1(n4826), .IN2(n5335), .IN3(n4958), .IN4(n2421), .IN5(
        g562), .IN6(n6110), .Q(g26895) );
  NOR2X0 U7189 ( .IN1(n4826), .IN2(n5335), .QN(n4958) );
  AO222X1 U7190 ( .IN1(n2982), .IN2(n5476), .IN3(n3273), .IN4(n2421), .IN5(
        g590), .IN6(n6097), .Q(g33538) );
  NOR2X0 U7191 ( .IN1(n2982), .IN2(n5476), .QN(n3273) );
  AO222X1 U7192 ( .IN1(n3745), .IN2(n5294), .IN3(n4200), .IN4(n2421), .IN5(
        g586), .IN6(n6108), .Q(g30334) );
  NOR2X0 U7193 ( .IN1(n3745), .IN2(n5294), .QN(n4200) );
  AO222X1 U7194 ( .IN1(n4201), .IN2(n5336), .IN3(n4536), .IN4(n2421), .IN5(
        g572), .IN6(n6105), .Q(g29224) );
  NOR2X0 U7195 ( .IN1(n4201), .IN2(n5336), .QN(n4536) );
  AO222X1 U7196 ( .IN1(n4537), .IN2(n5337), .IN3(n4825), .IN4(n2421), .IN5(
        g568), .IN6(n6108), .Q(g28045) );
  NOR2X0 U7197 ( .IN1(n4537), .IN2(n5337), .QN(n4825) );
  AO222X1 U7198 ( .IN1(n3274), .IN2(n5472), .IN3(n3683), .IN4(n2421), .IN5(
        g582), .IN6(n6100), .Q(g32978) );
  NOR2X0 U7199 ( .IN1(n3274), .IN2(n5472), .QN(n3683) );
  NAND4X0 U7200 ( .IN1(g1345), .IN2(g1367), .IN3(n1573), .IN4(g1379), .QN(
        n4896) );
  INVX0 U7201 ( .IN(n5067), .QN(n1573) );
  NAND4X0 U7202 ( .IN1(g1002), .IN2(g1024), .IN3(n5094), .IN4(g1036), .QN(
        n4921) );
  XNOR2X1 U7203 ( .IN1(g1339), .IN2(n5319), .Q(n5067) );
  AO221X1 U7204 ( .IN1(n6162), .IN2(n4797), .IN3(g2724), .IN4(n6086), .IN5(
        n2787), .Q(g28060) );
  XOR2X1 U7205 ( .IN1(g2729), .IN2(n4064), .Q(n4797) );
  AO221X1 U7206 ( .IN1(n4374), .IN2(g2735), .IN3(g2729), .IN4(n4375), .IN5(
        n2787), .Q(g29256) );
  NAND2X0 U7207 ( .IN1(n4376), .IN2(n6147), .QN(n4375) );
  NOR2X0 U7208 ( .IN1(g2729), .IN2(n6070), .QN(n4374) );
  XNOR2X1 U7209 ( .IN1(g2735), .IN2(n4064), .Q(n4376) );
  AO221X1 U7210 ( .IN1(g2712), .IN2(n6088), .IN3(n6177), .IN4(n5299), .IN5(
        n2787), .Q(g24263) );
  AO221X1 U7211 ( .IN1(n3095), .IN2(g2759), .IN3(test_so30), .IN4(n3096), 
        .IN5(n2787), .Q(g33608) );
  NAND2X0 U7212 ( .IN1(n3097), .IN2(n6149), .QN(n3096) );
  NOR2X0 U7213 ( .IN1(test_so30), .IN2(n6066), .QN(n3095) );
  XNOR2X1 U7214 ( .IN1(g2759), .IN2(n2790), .Q(n3097) );
  AO221X1 U7215 ( .IN1(n2785), .IN2(g2763), .IN3(g2759), .IN4(n2786), .IN5(
        n2787), .Q(g34022) );
  NAND2X0 U7216 ( .IN1(n2788), .IN2(n6180), .QN(n2786) );
  NOR2X0 U7217 ( .IN1(g2759), .IN2(n6063), .QN(n2785) );
  XOR2X1 U7218 ( .IN1(n2789), .IN2(g2763), .Q(n2788) );
  AO221X1 U7219 ( .IN1(n6157), .IN2(n3504), .IN3(g2748), .IN4(n6087), .IN5(
        n2787), .Q(g33019) );
  XNOR2X1 U7220 ( .IN1(n5300), .IN2(n2790), .Q(n3504) );
  XOR2X1 U7221 ( .IN1(g996), .IN2(n5320), .Q(n5094) );
  AO22X1 U7222 ( .IN1(g1536), .IN2(n6132), .IN3(n4164), .IN4(n1548), .Q(g30346) );
  NOR2X0 U7223 ( .IN1(n4165), .IN2(n6071), .QN(n4164) );
  XNOR2X1 U7224 ( .IN1(g1542), .IN2(n4166), .Q(n4165) );
  AO22X1 U7225 ( .IN1(g1193), .IN2(n6132), .IN3(n4182), .IN4(n1583), .Q(g30340) );
  NOR2X0 U7226 ( .IN1(n4183), .IN2(n6071), .QN(n4182) );
  XNOR2X1 U7227 ( .IN1(g1199), .IN2(n4184), .Q(n4183) );
  AO22X1 U7228 ( .IN1(g1542), .IN2(n6132), .IN3(n4161), .IN4(n1548), .Q(g30347) );
  NOR2X0 U7229 ( .IN1(n4162), .IN2(n6071), .QN(n4161) );
  XNOR2X1 U7230 ( .IN1(n4163), .IN2(g1413), .Q(n4162) );
  AO22X1 U7231 ( .IN1(g1199), .IN2(n6132), .IN3(n4179), .IN4(n1583), .Q(g30341) );
  NOR2X0 U7232 ( .IN1(n4180), .IN2(n6071), .QN(n4179) );
  XNOR2X1 U7233 ( .IN1(n4181), .IN2(g1070), .Q(n4180) );
  AO22X1 U7234 ( .IN1(g1514), .IN2(n4167), .IN3(n6337), .IN4(n4168), .Q(g30345) );
  NAND2X0 U7235 ( .IN1(n4170), .IN2(n6151), .QN(n4167) );
  NAND2X0 U7236 ( .IN1(n1548), .IN2(n3155), .QN(n4168) );
  XNOR2X1 U7237 ( .IN1(test_so49), .IN2(n6024), .Q(n4170) );
  AO22X1 U7238 ( .IN1(g1171), .IN2(n4185), .IN3(n6328), .IN4(n4186), .Q(g30339) );
  NAND2X0 U7239 ( .IN1(n4188), .IN2(n6170), .QN(n4185) );
  NAND2X0 U7240 ( .IN1(n1583), .IN2(n3235), .QN(n4186) );
  XNOR2X1 U7241 ( .IN1(g1183), .IN2(n6021), .Q(n4188) );
  AO22X1 U7242 ( .IN1(g1189), .IN2(n6128), .IN3(n6345), .IN4(n4917), .Q(g26918) );
  AO21X1 U7243 ( .IN1(g1193), .IN2(n4918), .IN3(n4191), .Q(n4917) );
  NAND2X0 U7244 ( .IN1(n4181), .IN2(g1070), .QN(n4918) );
  AO22X1 U7245 ( .IN1(g1532), .IN2(n6129), .IN3(n6342), .IN4(n4892), .Q(g26925) );
  AO21X1 U7246 ( .IN1(g1536), .IN2(n4893), .IN3(n4173), .Q(n4892) );
  NAND2X0 U7247 ( .IN1(n4163), .IN2(g1413), .QN(n4893) );
  ISOLANDX1 U7248 ( .D(n4172), .ISO(g1536), .Q(n4173) );
  ISOLANDX1 U7249 ( .D(n4190), .ISO(g1193), .Q(n4191) );
  AO22X1 U7250 ( .IN1(n6135), .IN2(g4388), .IN3(n4875), .IN4(n6294), .Q(g26947) );
  AO21X1 U7251 ( .IN1(n4872), .IN2(n4876), .IN3(n4871), .Q(n4875) );
  XNOR2X1 U7252 ( .IN1(g4375), .IN2(n5714), .Q(n4876) );
  AO21X1 U7253 ( .IN1(g4417), .IN2(n6122), .IN3(n4859), .Q(g26950) );
  AO21X1 U7254 ( .IN1(g4455), .IN2(n6122), .IN3(n4859), .Q(g26958) );
  NOR3X0 U7255 ( .IN1(g4392), .IN2(g4417), .IN3(n4872), .QN(n4871) );
  NOR2X0 U7256 ( .IN1(n5068), .IN2(n6079), .QN(g25631) );
  OA22X1 U7257 ( .IN1(n1837), .IN2(n5069), .IN3(n1574), .IN4(n5466), .Q(n5068)
         );
  OA221X1 U7258 ( .IN1(g1351), .IN2(n4896), .IN3(n5322), .IN4(n5070), .IN5(
        n4802), .Q(n5069) );
  OR2X1 U7259 ( .IN1(n5066), .IN2(g1389), .Q(n5070) );
  NOR2X0 U7260 ( .IN1(n5091), .IN2(n6079), .QN(g25622) );
  OA22X1 U7261 ( .IN1(n1927), .IN2(n5092), .IN3(n1928), .IN4(n5467), .Q(n5091)
         );
  OA221X1 U7262 ( .IN1(g1008), .IN2(n4921), .IN3(n5321), .IN4(n5093), .IN5(
        n4809), .Q(n5092) );
  OR2X1 U7263 ( .IN1(n5090), .IN2(g1046), .Q(n5093) );
  NAND2X0 U7264 ( .IN1(g2715), .IN2(n5465), .QN(n4411) );
  OR2X1 U7265 ( .IN1(n3557), .IN2(n5967), .Q(n3559) );
  AND3X1 U7266 ( .IN1(n3561), .IN2(n5511), .IN3(n3555), .Q(n5967) );
  NAND4X0 U7267 ( .IN1(n3373), .IN2(n3374), .IN3(n3375), .IN4(n3376), .QN(
        g34979) );
  OA22X1 U7268 ( .IN1(n3321), .IN2(DFF_420_n1), .IN3(n3364), .IN4(n5638), .Q(
        n3373) );
  OA22X1 U7269 ( .IN1(n3363), .IN2(n5981), .IN3(n3317), .IN4(n5308), .Q(n3375)
         );
  OA222X1 U7270 ( .IN1(n3345), .IN2(n5415), .IN3(n3320), .IN4(n5275), .IN5(
        n3344), .IN6(n5635), .Q(n3374) );
  NAND4X0 U7271 ( .IN1(n3329), .IN2(n3330), .IN3(n3331), .IN4(n3332), .QN(
        g34975) );
  OA22X1 U7272 ( .IN1(n3320), .IN2(n5643), .IN3(n3321), .IN4(DFF_829_n1), .Q(
        n3329) );
  OA222X1 U7273 ( .IN1(n3317), .IN2(n5495), .IN3(n3318), .IN4(n5344), .IN5(
        n3319), .IN6(n5295), .Q(n3330) );
  OA22X1 U7274 ( .IN1(n3334), .IN2(n6026), .IN3(n3335), .IN4(n6026), .Q(n3331)
         );
  NAND4X0 U7275 ( .IN1(n3353), .IN2(n3354), .IN3(n3355), .IN4(n3356), .QN(
        g34977) );
  OA22X1 U7276 ( .IN1(n3321), .IN2(DFF_1322_n1), .IN3(n3364), .IN4(n5639), .Q(
        n3353) );
  OA22X1 U7277 ( .IN1(g4737), .IN2(n3318), .IN3(g4927), .IN4(n3319), .Q(n3355)
         );
  OA222X1 U7278 ( .IN1(n3345), .IN2(n5286), .IN3(n3363), .IN4(n5493), .IN5(
        n3344), .IN6(n2549), .Q(n3354) );
  NAND4X0 U7279 ( .IN1(n5287), .IN2(n5327), .IN3(n5481), .IN4(n5109), .QN(
        n4955) );
  NOR3X0 U7280 ( .IN1(n4824), .IN2(g490), .IN3(g482), .QN(n5109) );
  OR2X1 U7281 ( .IN1(n3538), .IN2(n5968), .Q(n3540) );
  AND3X1 U7282 ( .IN1(n3542), .IN2(n5509), .IN3(n3536), .Q(n5968) );
  OR2X1 U7283 ( .IN1(n3595), .IN2(n5969), .Q(n3597) );
  AND3X1 U7284 ( .IN1(n3599), .IN2(n5507), .IN3(n3593), .Q(n5969) );
  OR2X1 U7285 ( .IN1(n3576), .IN2(n5970), .Q(n3578) );
  AND3X1 U7286 ( .IN1(n3580), .IN2(n5512), .IN3(n3574), .Q(n5970) );
  OR2X1 U7287 ( .IN1(n3613), .IN2(n5971), .Q(n3615) );
  AND3X1 U7288 ( .IN1(n3617), .IN2(n5510), .IN3(n3611), .Q(n5971) );
  OR2X1 U7289 ( .IN1(n3519), .IN2(n5972), .Q(n3521) );
  AND3X1 U7290 ( .IN1(n3523), .IN2(n5508), .IN3(n3517), .Q(n5972) );
  NAND4X0 U7291 ( .IN1(n3300), .IN2(n3301), .IN3(n3302), .IN4(n3303), .QN(
        g34970) );
  OA22X1 U7292 ( .IN1(n3320), .IN2(n5644), .IN3(n3321), .IN4(DFF_514_n1), .Q(
        n3300) );
  OA22X1 U7293 ( .IN1(n3308), .IN2(n6026), .IN3(n3310), .IN4(n6026), .Q(n3302)
         );
  OA222X1 U7294 ( .IN1(n3317), .IN2(n5641), .IN3(n3318), .IN4(n5312), .IN5(
        n3319), .IN6(n5408), .Q(n3301) );
  NAND4X0 U7295 ( .IN1(n3384), .IN2(n3385), .IN3(n3386), .IN4(n3387), .QN(
        g34971) );
  OA22X1 U7296 ( .IN1(n3321), .IN2(DFF_206_n1), .IN3(n3364), .IN4(n5640), .Q(
        n3384) );
  OA22X1 U7297 ( .IN1(n3363), .IN2(n5983), .IN3(n3317), .IN4(n5377), .Q(n3386)
         );
  OA222X1 U7298 ( .IN1(n3345), .IN2(n5409), .IN3(n3320), .IN4(n5307), .IN5(
        n3344), .IN6(n5623), .Q(n3385) );
  NAND4X0 U7299 ( .IN1(n3365), .IN2(n3366), .IN3(n3367), .IN4(n3368), .QN(
        g34978) );
  OA22X1 U7300 ( .IN1(n3321), .IN2(DFF_1012_n1), .IN3(n3364), .IN4(n5484), .Q(
        n3365) );
  OA22X1 U7301 ( .IN1(n3363), .IN2(n5494), .IN3(n3317), .IN4(n5347), .Q(n3367)
         );
  OA222X1 U7302 ( .IN1(g952), .IN2(n3345), .IN3(n3320), .IN4(n5487), .IN5(
        g1296), .IN6(n3344), .Q(n3366) );
  NAND4X0 U7303 ( .IN1(n3322), .IN2(n3323), .IN3(n3324), .IN4(n3325), .QN(
        g34974) );
  OA22X1 U7304 ( .IN1(n3320), .IN2(n5499), .IN3(n3321), .IN4(DFF_477_n1), .Q(
        n3322) );
  OA222X1 U7305 ( .IN1(n3317), .IN2(n5496), .IN3(n3318), .IN4(n5296), .IN5(
        n3319), .IN6(n5346), .Q(n3323) );
  OA22X1 U7306 ( .IN1(n3326), .IN2(n6026), .IN3(n3327), .IN4(n6026), .Q(n3324)
         );
  NAND4X0 U7307 ( .IN1(n3340), .IN2(n3341), .IN3(n3342), .IN4(n3343), .QN(
        g34976) );
  OA22X1 U7308 ( .IN1(n3320), .IN2(n5498), .IN3(n3321), .IN4(DFF_150_n1), .Q(
        n3340) );
  OA22X1 U7309 ( .IN1(n3346), .IN2(n6026), .IN3(n3347), .IN4(n6026), .Q(n3342)
         );
  OA222X1 U7310 ( .IN1(n3317), .IN2(n5497), .IN3(n3318), .IN4(n5345), .IN5(
        n3319), .IN6(n5297), .Q(n3341) );
  XNOR3X1 U7311 ( .IN1(n2399), .IN2(n2400), .IN3(n2401), .Q(n2393) );
  OA21X1 U7312 ( .IN1(g24163), .IN2(n5954), .IN3(g55), .Q(n2399) );
  XNOR3X1 U7313 ( .IN1(n2402), .IN2(g34979), .IN3(g34971), .Q(n2401) );
  XNOR3X1 U7314 ( .IN1(g34970), .IN2(n1456), .IN3(n2403), .Q(n2400) );
  NAND2X0 U7315 ( .IN1(g22), .IN2(n2393), .QN(g34972) );
  NAND2X0 U7316 ( .IN1(g22), .IN2(n1309), .QN(g34927) );
  NAND2X0 U7317 ( .IN1(g22), .IN2(n1452), .QN(g34925) );
  NAND2X0 U7318 ( .IN1(g22), .IN2(n1453), .QN(g34923) );
  NAND2X0 U7319 ( .IN1(g22), .IN2(n1454), .QN(g34921) );
  NAND2X0 U7320 ( .IN1(g22), .IN2(n1455), .QN(g34919) );
  NAND2X0 U7321 ( .IN1(g22), .IN2(n1456), .QN(g34917) );
  NAND2X0 U7322 ( .IN1(g22), .IN2(n1277), .QN(g34915) );
  NAND2X0 U7323 ( .IN1(g22), .IN2(n1457), .QN(g34913) );
  OA21X1 U7324 ( .IN1(g3845), .IN2(g3831), .IN3(n6353), .Q(n4853) );
  XNOR2X1 U7325 ( .IN1(g4322), .IN2(n5962), .Q(n3094) );
  NAND2X0 U7326 ( .IN1(g376), .IN2(g358), .QN(n5125) );
  NOR2X0 U7327 ( .IN1(n6082), .IN2(g4392), .QN(n4863) );
  AND3X1 U7328 ( .IN1(n1489), .IN2(g4311), .IN3(n3060), .Q(n2761) );
  NAND2X0 U7329 ( .IN1(g5124), .IN2(n6164), .QN(n3764) );
  AND3X1 U7330 ( .IN1(g4849), .IN2(g4843), .IN3(g4859), .Q(n3013) );
  AND3X1 U7331 ( .IN1(g4659), .IN2(test_so19), .IN3(g4669), .Q(n3012) );
  AND3X1 U7332 ( .IN1(test_so60), .IN2(n4198), .IN3(n4199), .Q(n3743) );
  NAND2X0 U7333 ( .IN1(g385), .IN2(n2077), .QN(n5121) );
  AO21X1 U7334 ( .IN1(g2886), .IN2(n6120), .IN3(n2460), .Q(g34800) );
  NAND2X0 U7335 ( .IN1(n1802), .IN2(g34979), .QN(n2461) );
  NAND3X0 U7336 ( .IN1(g4776), .IN2(n5285), .IN3(g4793), .QN(n4314) );
  NAND3X0 U7337 ( .IN1(g4966), .IN2(n5284), .IN3(g4983), .QN(n4292) );
  NAND4X0 U7338 ( .IN1(n1539), .IN2(n4831), .IN3(n4832), .IN4(n4833), .QN(
        n4205) );
  NAND2X0 U7339 ( .IN1(g807), .IN2(g554), .QN(n4831) );
  OR3X1 U7340 ( .IN1(g718), .IN2(g753), .IN3(g655), .Q(n4832) );
  NAND3X0 U7341 ( .IN1(g718), .IN2(g655), .IN3(g753), .QN(n4833) );
  OA221X1 U7342 ( .IN1(n3369), .IN2(n6026), .IN3(n3370), .IN4(n6026), .IN5(
        n3333), .Q(n3368) );
  OA221X1 U7343 ( .IN1(g550), .IN2(n3311), .IN3(n3312), .IN4(n5471), .IN5(
        n3372), .Q(n3369) );
  OA221X1 U7344 ( .IN1(n2545), .IN2(n5342), .IN3(n3337), .IN4(n5488), .IN5(
        n3371), .Q(n3370) );
  OA222X1 U7345 ( .IN1(n3352), .IN2(n5292), .IN3(n3314), .IN4(n5337), .IN5(
        n3315), .IN6(n5475), .Q(n3372) );
  OA221X1 U7346 ( .IN1(n3377), .IN2(n6026), .IN3(n3378), .IN4(n6025), .IN5(
        n3333), .Q(n3376) );
  NOR2X0 U7347 ( .IN1(n3379), .IN2(n3380), .QN(n3378) );
  OA221X1 U7348 ( .IN1(g30329), .IN2(n3311), .IN3(n3312), .IN4(n5470), .IN5(
        n3383), .Q(n3377) );
  AO222X1 U7349 ( .IN1(g24182), .IN2(n1800), .IN3(test_so14), .IN4(n1802), 
        .IN5(g24171), .IN6(n1801), .Q(n3380) );
  OA221X1 U7350 ( .IN1(n3357), .IN2(n6026), .IN3(n3358), .IN4(n6026), .IN5(
        n3333), .Q(n3356) );
  NOR2X0 U7351 ( .IN1(n3360), .IN2(n3361), .QN(n3357) );
  OA221X1 U7352 ( .IN1(n3311), .IN2(n5490), .IN3(n3312), .IN4(n5331), .IN5(
        n3359), .Q(n3358) );
  AO222X1 U7353 ( .IN1(g2868), .IN2(n1800), .IN3(g2882), .IN4(n1793), .IN5(
        n1801), .IN6(g37), .Q(n3361) );
  INVX0 U7354 ( .IN(n6684), .QN(n6678) );
  INVX0 U7355 ( .IN(g35), .QN(n6684) );
  INVX0 U7356 ( .IN(g35), .QN(n6682) );
  AO221X1 U7357 ( .IN1(g1624), .IN2(n3649), .IN3(n1398), .IN4(test_so94), 
        .IN5(n3648), .Q(g32988) );
  AO221X1 U7358 ( .IN1(g2028), .IN2(n3596), .IN3(n1395), .IN4(g2051), .IN5(
        n3595), .Q(g33000) );
  AO221X1 U7359 ( .IN1(g1760), .IN2(n3631), .IN3(n1397), .IN4(g1783), .IN5(
        n3630), .Q(g32992) );
  AO221X1 U7360 ( .IN1(g2185), .IN2(n3577), .IN3(n1394), .IN4(g2208), .IN5(
        n3576), .Q(g33004) );
  AO221X1 U7361 ( .IN1(g2453), .IN2(n3539), .IN3(n1392), .IN4(g2476), .IN5(
        n3538), .Q(g33012) );
  AO221X1 U7362 ( .IN1(g2319), .IN2(n3558), .IN3(n1393), .IN4(test_so21), 
        .IN5(n3557), .Q(g33008) );
  AO221X1 U7363 ( .IN1(g2587), .IN2(n3520), .IN3(n1391), .IN4(g2610), .IN5(
        n3519), .Q(g33016) );
  AO221X1 U7364 ( .IN1(g1894), .IN2(n3614), .IN3(n1396), .IN4(g1917), .IN5(
        n3613), .Q(g32996) );
  AO21X1 U7365 ( .IN1(g4297), .IN2(n6121), .IN3(n2488), .Q(g34735) );
  AO21X1 U7366 ( .IN1(test_so41), .IN2(n6121), .IN3(n2510), .Q(g34723) );
  AO21X1 U7367 ( .IN1(g2848), .IN2(n6121), .IN3(n2480), .Q(g34793) );
  OR2X1 U7368 ( .IN1(n2440), .IN2(g2856), .Q(n2481) );
  AO21X1 U7369 ( .IN1(g2873), .IN2(n6120), .IN3(n2462), .Q(g34799) );
  AO21X1 U7370 ( .IN1(g4172), .IN2(n6121), .IN3(n2490), .Q(g34734) );
  AO21X1 U7371 ( .IN1(g2902), .IN2(n6120), .IN3(n2452), .Q(g34802) );
  OR2X1 U7372 ( .IN1(n2455), .IN2(g2917), .Q(n2454) );
  AO21X1 U7373 ( .IN1(g534), .IN2(n6121), .IN3(n2514), .Q(g34720) );
  AO21X1 U7374 ( .IN1(g2898), .IN2(n6121), .IN3(n2466), .Q(g34796) );
  OR2X1 U7375 ( .IN1(n2433), .IN2(g2882), .Q(n2467) );
  AO21X1 U7376 ( .IN1(g2882), .IN2(n6120), .IN3(n2465), .Q(g34797) );
  AO21X1 U7377 ( .IN1(g21292), .IN2(n6122), .IN3(n2513), .Q(g34721) );
  AO21X1 U7378 ( .IN1(g2970), .IN2(n6119), .IN3(n2456), .Q(g34801) );
  OR2X1 U7379 ( .IN1(g2902), .IN2(g301), .Q(n2458) );
  AO21X1 U7380 ( .IN1(g2965), .IN2(n6120), .IN3(n2446), .Q(g34804) );
  NAND2X0 U7381 ( .IN1(n2449), .IN2(n5750), .QN(n2448) );
  AO21X1 U7382 ( .IN1(g20652), .IN2(n6121), .IN3(n2482), .Q(g34792) );
  OR2X1 U7383 ( .IN1(n2442), .IN2(g2848), .Q(n2483) );
  AO21X1 U7384 ( .IN1(g1296), .IN2(n6119), .IN3(n2497), .Q(g34730) );
  AO21X1 U7385 ( .IN1(g2878), .IN2(n6121), .IN3(n2463), .Q(g34798) );
  AO21X1 U7386 ( .IN1(g2864), .IN2(n6120), .IN3(n2468), .Q(g34795) );
  AO21X1 U7387 ( .IN1(g2927), .IN2(n6120), .IN3(n2443), .Q(g34806) );
  OR2X1 U7388 ( .IN1(g4072), .IN2(g4153), .Q(n2444) );
  AO21X1 U7389 ( .IN1(g952), .IN2(n6121), .IN3(n2503), .Q(g34727) );
  AO21X1 U7390 ( .IN1(g2941), .IN2(n6120), .IN3(n2434), .Q(g34807) );
  OR4X1 U7391 ( .IN1(n2441), .IN2(n2442), .IN3(g2946), .IN4(g2955), .Q(n2435)
         );
  OR4X1 U7392 ( .IN1(n2437), .IN2(n2438), .IN3(n2439), .IN4(n2440), .Q(n2436)
         );
  OA21X1 U7393 ( .IN1(g6537), .IN2(g6523), .IN3(n6357), .Q(n4849) );
  AO222X1 U7394 ( .IN1(n4015), .IN2(n1732), .IN3(n4019), .IN4(g3251), .IN5(
        g3235), .IN6(n6114), .Q(g30407) );
  OA21X1 U7395 ( .IN1(n4020), .IN2(n3500), .IN3(n6374), .Q(n4019) );
  AO222X1 U7396 ( .IN1(n3908), .IN2(n1576), .IN3(n3912), .IN4(g5260), .IN5(
        g5244), .IN6(n6095), .Q(g30473) );
  OA21X1 U7397 ( .IN1(n3904), .IN2(n3444), .IN3(n6386), .Q(n3912) );
  AO222X1 U7398 ( .IN1(n4027), .IN2(n1729), .IN3(n4029), .IN4(g3223), .IN5(
        g3199), .IN6(n6114), .Q(g30400) );
  OA21X1 U7399 ( .IN1(n3501), .IN2(n3495), .IN3(n6383), .Q(n4029) );
  AO222X1 U7400 ( .IN1(n4037), .IN2(n6038), .IN3(n4038), .IN4(g3191), .IN5(
        test_so88), .IN6(n6115), .Q(g30395) );
  NOR2X0 U7401 ( .IN1(n4037), .IN2(n6073), .QN(n4038) );
  ISOLANDX1 U7402 ( .D(n4034), .ISO(n4020), .Q(n4037) );
  AO222X1 U7403 ( .IN1(n4039), .IN2(n6029), .IN3(n4040), .IN4(g3187), .IN5(
        g3179), .IN6(n6114), .Q(g30394) );
  NOR2X0 U7404 ( .IN1(n4039), .IN2(n6073), .QN(n4040) );
  ISOLANDX1 U7405 ( .D(n4034), .ISO(n4014), .Q(n4039) );
  AO222X1 U7406 ( .IN1(n3808), .IN2(n1510), .IN3(n3813), .IN4(g6295), .IN5(
        g6279), .IN6(n6092), .Q(g30535) );
  OA21X1 U7407 ( .IN1(n3414), .IN2(n3807), .IN3(n6398), .Q(n3813) );
  AO222X1 U7408 ( .IN1(n4009), .IN2(n6033), .IN3(n4010), .IN4(g3211), .IN5(
        g3255), .IN6(n6113), .Q(g30412) );
  NOR2X0 U7409 ( .IN1(n4009), .IN2(n6074), .QN(n4010) );
  NOR2X0 U7410 ( .IN1(n3495), .IN2(n5652), .QN(n4009) );
  AO222X1 U7411 ( .IN1(n3972), .IN2(n6037), .IN3(n3973), .IN4(g3893), .IN5(
        g3897), .IN6(n6112), .Q(g30437) );
  NOR2X0 U7412 ( .IN1(n3972), .IN2(n6075), .QN(n3973) );
  ISOLANDX1 U7413 ( .D(n3969), .ISO(n3947), .Q(n3972) );
  AO222X1 U7414 ( .IN1(n3929), .IN2(n6040), .IN3(n3930), .IN4(g5200), .IN5(
        g5204), .IN6(n6113), .Q(g30461) );
  NOR2X0 U7415 ( .IN1(n3929), .IN2(n6066), .QN(n3930) );
  ISOLANDX1 U7416 ( .D(n3926), .ISO(n3904), .Q(n3929) );
  AO222X1 U7417 ( .IN1(n3951), .IN2(n1903), .IN3(n3955), .IN4(g3953), .IN5(
        g3937), .IN6(n6111), .Q(g30449) );
  OA21X1 U7418 ( .IN1(n3947), .IN2(n3479), .IN3(n6382), .Q(n3955) );
  AO222X1 U7419 ( .IN1(n3808), .IN2(n1509), .IN3(n3812), .IN4(g6299), .IN5(
        g6283), .IN6(n6105), .Q(g30536) );
  OA21X1 U7420 ( .IN1(n3804), .IN2(n3414), .IN3(n6398), .Q(n3812) );
  AO222X1 U7421 ( .IN1(n3881), .IN2(n1968), .IN3(n3882), .IN4(g5599), .IN5(
        g5583), .IN6(n6093), .Q(g30492) );
  OA21X1 U7422 ( .IN1(n3877), .IN2(n3436), .IN3(n6389), .Q(n3882) );
  AO222X1 U7423 ( .IN1(n3785), .IN2(n2222), .IN3(n3787), .IN4(g6617), .IN5(
        g6593), .IN6(n6103), .Q(g30550) );
  OA21X1 U7424 ( .IN1(n3768), .IN2(n3407), .IN3(n6400), .Q(n3787) );
  AO222X1 U7425 ( .IN1(n3863), .IN2(n6043), .IN3(n3864), .IN4(g5893), .IN5(
        g5897), .IN6(n6092), .Q(g30503) );
  NOR2X0 U7426 ( .IN1(n3863), .IN2(n6073), .QN(n3864) );
  ISOLANDX1 U7427 ( .D(n3860), .ISO(n3838), .Q(n3863) );
  AO222X1 U7428 ( .IN1(n4015), .IN2(n1729), .IN3(n4018), .IN4(g3255), .IN5(
        g3239), .IN6(n6114), .Q(g30408) );
  OA21X1 U7429 ( .IN1(n3500), .IN2(n3495), .IN3(n6374), .Q(n4018) );
  AO222X1 U7430 ( .IN1(n3943), .IN2(n6039), .IN3(n3944), .IN4(g3913), .IN5(
        g3957), .IN6(n6111), .Q(g30454) );
  NOR2X0 U7431 ( .IN1(n3943), .IN2(n6076), .QN(n3944) );
  NOR2X0 U7432 ( .IN1(n3945), .IN2(n5648), .QN(n3943) );
  AO222X1 U7433 ( .IN1(n4012), .IN2(n6038), .IN3(n4013), .IN4(test_so88), 
        .IN5(g3247), .IN6(n6114), .Q(g30410) );
  NOR2X0 U7434 ( .IN1(n4012), .IN2(n6073), .QN(n4013) );
  NOR2X0 U7435 ( .IN1(n4014), .IN2(n5652), .QN(n4012) );
  AO222X1 U7436 ( .IN1(n4003), .IN2(n6039), .IN3(n4004), .IN4(g3550), .IN5(
        g3554), .IN6(n6113), .Q(g30417) );
  NOR2X0 U7437 ( .IN1(n4003), .IN2(n6074), .QN(n4004) );
  ISOLANDX1 U7438 ( .D(n4002), .ISO(n3978), .Q(n4003) );
  AO222X1 U7439 ( .IN1(n3842), .IN2(n1816), .IN3(n3846), .IN4(g5953), .IN5(
        g5937), .IN6(n6090), .Q(g30515) );
  OA21X1 U7440 ( .IN1(n3838), .IN2(n3424), .IN3(n6394), .Q(n3846) );
  AO222X1 U7441 ( .IN1(n3990), .IN2(n1680), .IN3(n3991), .IN4(g3594), .IN5(
        g3578), .IN6(n6112), .Q(g30426) );
  OA21X1 U7442 ( .IN1(n3986), .IN2(n3491), .IN3(n6377), .Q(n3991) );
  AO222X1 U7443 ( .IN1(n4027), .IN2(n1731), .IN3(n4031), .IN4(g3215), .IN5(
        g3187), .IN6(n6115), .Q(g30398) );
  OA21X1 U7444 ( .IN1(n3501), .IN2(n4014), .IN3(n6404), .Q(n4031) );
  AO222X1 U7445 ( .IN1(n4015), .IN2(n1730), .IN3(n4016), .IN4(test_so84), 
        .IN5(g3243), .IN6(n6114), .Q(g30409) );
  OA21X1 U7446 ( .IN1(n4017), .IN2(n3500), .IN3(n6374), .Q(n4016) );
  AO222X1 U7447 ( .IN1(n4032), .IN2(n6031), .IN3(n4033), .IN4(g3207), .IN5(
        g3211), .IN6(n6114), .Q(g30397) );
  NOR2X0 U7448 ( .IN1(n4032), .IN2(n6073), .QN(n4033) );
  ISOLANDX1 U7449 ( .D(n4034), .ISO(n4017), .Q(n4032) );
  AO222X1 U7450 ( .IN1(n3834), .IN2(n6044), .IN3(n3835), .IN4(g5913), .IN5(
        g5957), .IN6(n6089), .Q(g30520) );
  NOR2X0 U7451 ( .IN1(n3834), .IN2(n6072), .QN(n3835) );
  NOR2X0 U7452 ( .IN1(n3836), .IN2(n5649), .QN(n3834) );
  AO222X1 U7453 ( .IN1(n4035), .IN2(n6030), .IN3(n4036), .IN4(g3199), .IN5(
        g3203), .IN6(n6114), .Q(g30396) );
  NOR2X0 U7454 ( .IN1(n4035), .IN2(n6073), .QN(n4036) );
  ISOLANDX1 U7455 ( .D(n4034), .ISO(n3495), .Q(n4035) );
  AO222X1 U7456 ( .IN1(n3919), .IN2(n1576), .IN3(n3922), .IN4(test_so82), 
        .IN5(g5200), .IN6(n6096), .Q(g30465) );
  OA21X1 U7457 ( .IN1(n3904), .IN2(n3447), .IN3(n6383), .Q(n3922) );
  AO222X1 U7458 ( .IN1(n3984), .IN2(n1680), .IN3(n3985), .IN4(g3610), .IN5(
        g3594), .IN6(n6112), .Q(g30430) );
  OA21X1 U7459 ( .IN1(n3986), .IN2(n3489), .IN3(n6378), .Q(n3985) );
  AO222X1 U7460 ( .IN1(n3400), .IN2(n6046), .IN3(n3769), .IN4(g6597), .IN5(
        g6645), .IN6(n6102), .Q(g30561) );
  NOR2X0 U7461 ( .IN1(n3400), .IN2(n6070), .QN(n3769) );
  AO222X1 U7462 ( .IN1(n3797), .IN2(n6045), .IN3(n3798), .IN4(g6581), .IN5(
        g6573), .IN6(n6104), .Q(g30544) );
  NOR2X0 U7463 ( .IN1(n3797), .IN2(n6071), .QN(n3798) );
  ISOLANDX1 U7464 ( .D(n3792), .ISO(n3773), .Q(n3797) );
  AO222X1 U7465 ( .IN1(n3790), .IN2(n6045), .IN3(n3791), .IN4(g6601), .IN5(
        g6605), .IN6(n6104), .Q(g30547) );
  NOR2X0 U7466 ( .IN1(n3790), .IN2(n6071), .QN(n3791) );
  ISOLANDX1 U7467 ( .D(n3792), .ISO(n3776), .Q(n3790) );
  AO222X1 U7468 ( .IN1(n4027), .IN2(n1732), .IN3(n4030), .IN4(g3219), .IN5(
        g3191), .IN6(n6115), .Q(g30399) );
  OA21X1 U7469 ( .IN1(n4020), .IN2(n3501), .IN3(n6403), .Q(n4030) );
  AO222X1 U7470 ( .IN1(n3962), .IN2(n1903), .IN3(n3965), .IN4(g3921), .IN5(
        g3893), .IN6(n6111), .Q(g30441) );
  OA21X1 U7471 ( .IN1(n3947), .IN2(n3482), .IN3(n6379), .Q(n3965) );
  AO222X1 U7472 ( .IN1(n3808), .IN2(n1511), .IN3(n3811), .IN4(g6303), .IN5(
        g6287), .IN6(n6105), .Q(g30537) );
  OA21X1 U7473 ( .IN1(n3802), .IN2(n3414), .IN3(n6399), .Q(n3811) );
  AO222X1 U7474 ( .IN1(n3914), .IN2(n1581), .IN3(n3915), .IN4(g5252), .IN5(
        g5236), .IN6(n6096), .Q(g30471) );
  OA21X1 U7475 ( .IN1(n3910), .IN2(n3446), .IN3(n6385), .Q(n3915) );
  AO222X1 U7476 ( .IN1(n3853), .IN2(n1816), .IN3(n3856), .IN4(g5921), .IN5(
        g5893), .IN6(n6091), .Q(g30507) );
  OA21X1 U7477 ( .IN1(n3838), .IN2(n3427), .IN3(n6391), .Q(n3856) );
  AO222X1 U7478 ( .IN1(n3440), .IN2(n6041), .IN3(n3903), .IN4(g5212), .IN5(
        g5260), .IN6(n6095), .Q(g30477) );
  NOR2X0 U7479 ( .IN1(n3440), .IN2(n6076), .QN(n3903) );
  AO222X1 U7480 ( .IN1(n3795), .IN2(n6045), .IN3(n3796), .IN4(test_so71), 
        .IN5(g6589), .IN6(n6104), .Q(g30545) );
  NOR2X0 U7481 ( .IN1(n3795), .IN2(n6071), .QN(n3796) );
  ISOLANDX1 U7482 ( .D(n3792), .ISO(n3770), .Q(n3795) );
  AO222X1 U7483 ( .IN1(n3766), .IN2(n6037), .IN3(n3767), .IN4(g6605), .IN5(
        g6649), .IN6(n6102), .Q(g30562) );
  NOR2X0 U7484 ( .IN1(n3766), .IN2(n6070), .QN(n3767) );
  NOR2X0 U7485 ( .IN1(n3768), .IN2(n5646), .QN(n3766) );
  AO222X1 U7486 ( .IN1(n3957), .IN2(n1908), .IN3(n3958), .IN4(g3945), .IN5(
        g3929), .IN6(n6111), .Q(g30447) );
  OA21X1 U7487 ( .IN1(n3953), .IN2(n3481), .IN3(n6381), .Q(n3958) );
  AO222X1 U7488 ( .IN1(n3819), .IN2(n1510), .IN3(n3823), .IN4(g6263), .IN5(
        g6235), .IN6(n6089), .Q(g30527) );
  OA21X1 U7489 ( .IN1(n3807), .IN2(n3417), .IN3(n6395), .Q(n3823) );
  AO222X1 U7490 ( .IN1(n3891), .IN2(n6042), .IN3(n3892), .IN4(g5563), .IN5(
        g5567), .IN6(n6094), .Q(g30484) );
  NOR2X0 U7491 ( .IN1(n3891), .IN2(n6074), .QN(n3892) );
  ISOLANDX1 U7492 ( .D(n3893), .ISO(n3877), .Q(n3891) );
  AO222X1 U7493 ( .IN1(n3962), .IN2(n1905), .IN3(n3964), .IN4(g3925), .IN5(
        g3901), .IN6(n6111), .Q(g30442) );
  OA21X1 U7494 ( .IN1(n3945), .IN2(n3482), .IN3(n6379), .Q(n3964) );
  AO222X1 U7495 ( .IN1(n3919), .IN2(n1581), .IN3(n3920), .IN4(g5236), .IN5(
        g5216), .IN6(n6096), .Q(g30467) );
  OA21X1 U7496 ( .IN1(n3910), .IN2(n3447), .IN3(n6384), .Q(n3920) );
  AO222X1 U7497 ( .IN1(n3981), .IN2(n6036), .IN3(n3982), .IN4(g3546), .IN5(
        g3598), .IN6(n6112), .Q(g30431) );
  NOR2X0 U7498 ( .IN1(n3981), .IN2(n6075), .QN(n3982) );
  NOR2X0 U7499 ( .IN1(n3983), .IN2(n5645), .QN(n3981) );
  AO222X1 U7500 ( .IN1(n3771), .IN2(n6046), .IN3(n3772), .IN4(g6589), .IN5(
        g6641), .IN6(n6103), .Q(g30560) );
  NOR2X0 U7501 ( .IN1(n3771), .IN2(n6070), .QN(n3772) );
  NOR2X0 U7502 ( .IN1(n3773), .IN2(n5646), .QN(n3771) );
  AO222X1 U7503 ( .IN1(n3785), .IN2(n2225), .IN3(n3789), .IN4(g6609), .IN5(
        g6581), .IN6(n6104), .Q(g30548) );
  OA21X1 U7504 ( .IN1(n3773), .IN2(n3407), .IN3(n6400), .Q(n3789) );
  AO222X1 U7505 ( .IN1(n3914), .IN2(n1576), .IN3(n3917), .IN4(g5244), .IN5(
        test_so82), .IN6(n6096), .Q(g30469) );
  OA21X1 U7506 ( .IN1(n3904), .IN2(n3446), .IN3(n6385), .Q(n3917) );
  AO222X1 U7507 ( .IN1(n3848), .IN2(n1821), .IN3(n3849), .IN4(g5945), .IN5(
        g5929), .IN6(n6090), .Q(g30513) );
  OA21X1 U7508 ( .IN1(n3844), .IN2(n3426), .IN3(n6393), .Q(n3849) );
  AO222X1 U7509 ( .IN1(n3951), .IN2(n1904), .IN3(n3956), .IN4(test_so65), 
        .IN5(g3933), .IN6(n6111), .Q(g30448) );
  OA21X1 U7510 ( .IN1(n3479), .IN2(n3950), .IN3(n6381), .Q(n3956) );
  AO222X1 U7511 ( .IN1(n3827), .IN2(n6044), .IN3(n3828), .IN4(g6247), .IN5(
        g6251), .IN6(n6089), .Q(g30525) );
  NOR2X0 U7512 ( .IN1(n3827), .IN2(n6072), .QN(n3828) );
  ISOLANDX1 U7513 ( .D(n3826), .ISO(n3802), .Q(n3827) );
  AO222X1 U7514 ( .IN1(n3896), .IN2(n6041), .IN3(n3897), .IN4(g5547), .IN5(
        g5551), .IN6(n6094), .Q(g30482) );
  NOR2X0 U7515 ( .IN1(n3896), .IN2(n6075), .QN(n3897) );
  ISOLANDX1 U7516 ( .D(n3893), .ISO(n3871), .Q(n3896) );
  AO222X1 U7517 ( .IN1(n3919), .IN2(n1577), .IN3(n3923), .IN4(g5224), .IN5(
        g5196), .IN6(n6096), .Q(g30464) );
  OA21X1 U7518 ( .IN1(n3907), .IN2(n3447), .IN3(n6383), .Q(n3923) );
  AO222X1 U7519 ( .IN1(n3853), .IN2(n1818), .IN3(n3855), .IN4(g5925), .IN5(
        g5901), .IN6(n6091), .Q(g30508) );
  OA21X1 U7520 ( .IN1(n3836), .IN2(n3427), .IN3(n6392), .Q(n3855) );
  AO222X1 U7521 ( .IN1(n3962), .IN2(n1908), .IN3(n3963), .IN4(g3929), .IN5(
        g3909), .IN6(n6111), .Q(g30443) );
  OA21X1 U7522 ( .IN1(n3953), .IN2(n3482), .IN3(n6380), .Q(n3963) );
  AO222X1 U7523 ( .IN1(n3814), .IN2(n1509), .IN3(n3817), .IN4(g6283), .IN5(
        g6267), .IN6(n6089), .Q(g30532) );
  OA21X1 U7524 ( .IN1(n3804), .IN2(n3416), .IN3(n6397), .Q(n3817) );
  AO222X1 U7525 ( .IN1(n3886), .IN2(n1968), .IN3(n3887), .IN4(g5583), .IN5(
        g5563), .IN6(n6093), .Q(g30488) );
  OA21X1 U7526 ( .IN1(n3877), .IN2(n3437), .IN3(n6388), .Q(n3887) );
  AO222X1 U7527 ( .IN1(n3875), .IN2(n1969), .IN3(n3880), .IN4(g5603), .IN5(
        g5587), .IN6(n6093), .Q(g30493) );
  OA21X1 U7528 ( .IN1(n3434), .IN2(n3874), .IN3(n6390), .Q(n3880) );
  AO222X1 U7529 ( .IN1(n3842), .IN2(n1817), .IN3(n3847), .IN4(g5949), .IN5(
        g5933), .IN6(n6090), .Q(g30514) );
  OA21X1 U7530 ( .IN1(n3424), .IN2(n3841), .IN3(n6394), .Q(n3847) );
  AO222X1 U7531 ( .IN1(n3957), .IN2(n1903), .IN3(n3960), .IN4(g3937), .IN5(
        g3921), .IN6(n6111), .Q(g30445) );
  OA21X1 U7532 ( .IN1(n3947), .IN2(n3481), .IN3(n6380), .Q(n3960) );
  AO222X1 U7533 ( .IN1(n3853), .IN2(n1821), .IN3(n3854), .IN4(g5929), .IN5(
        g5909), .IN6(n6091), .Q(g30509) );
  OA21X1 U7534 ( .IN1(n3844), .IN2(n3427), .IN3(n6392), .Q(n3854) );
  AO222X1 U7535 ( .IN1(n3848), .IN2(n1816), .IN3(n3851), .IN4(g5937), .IN5(
        g5921), .IN6(n6091), .Q(g30511) );
  OA21X1 U7536 ( .IN1(n3838), .IN2(n3426), .IN3(n6393), .Q(n3851) );
  AO222X1 U7537 ( .IN1(n3774), .IN2(n2224), .IN3(n3775), .IN4(g6653), .IN5(
        g6637), .IN6(n6103), .Q(g30559) );
  OA21X1 U7538 ( .IN1(n3776), .IN2(n3404), .IN3(n6403), .Q(n3775) );
  AO222X1 U7539 ( .IN1(n3900), .IN2(n6041), .IN3(n3901), .IN4(g5220), .IN5(
        g5264), .IN6(n6095), .Q(g30478) );
  NOR2X0 U7540 ( .IN1(n3900), .IN2(n6075), .QN(n3901) );
  NOR2X0 U7541 ( .IN1(n3902), .IN2(n5650), .QN(n3900) );
  AO222X1 U7542 ( .IN1(n3976), .IN2(n6037), .IN3(n3977), .IN4(g3562), .IN5(
        g3606), .IN6(n6112), .Q(g30433) );
  NOR2X0 U7543 ( .IN1(n3976), .IN2(n6075), .QN(n3977) );
  NOR2X0 U7544 ( .IN1(n3978), .IN2(n5645), .QN(n3976) );
  AO222X1 U7545 ( .IN1(n3785), .IN2(n2226), .IN3(n3788), .IN4(g6613), .IN5(
        test_so71), .IN6(n6103), .Q(g30549) );
  OA21X1 U7546 ( .IN1(n3770), .IN2(n3407), .IN3(n6399), .Q(n3788) );
  AO222X1 U7547 ( .IN1(n4007), .IN2(n6034), .IN3(n4008), .IN4(g3538), .IN5(
        g3530), .IN6(n6113), .Q(g30415) );
  NOR2X0 U7548 ( .IN1(n4007), .IN2(n6074), .QN(n4008) );
  ISOLANDX1 U7549 ( .D(n4002), .ISO(n3983), .Q(n4007) );
  AO222X1 U7550 ( .IN1(n4015), .IN2(n1731), .IN3(n4021), .IN4(g3247), .IN5(
        g3231), .IN6(n6115), .Q(g30406) );
  OA21X1 U7551 ( .IN1(n3500), .IN2(n4014), .IN3(n6373), .Q(n4021) );
  AO222X1 U7552 ( .IN1(n3908), .IN2(n1577), .IN3(n3913), .IN4(g5256), .IN5(
        g5240), .IN6(n6095), .Q(g30472) );
  OA21X1 U7553 ( .IN1(n3444), .IN2(n3907), .IN3(n6386), .Q(n3913) );
  AO222X1 U7554 ( .IN1(n1544), .IN2(n6032), .IN3(n4011), .IN4(g3203), .IN5(
        g3251), .IN6(n6114), .Q(g30411) );
  NOR2X0 U7555 ( .IN1(n1544), .IN2(n6074), .QN(n4011) );
  INVX0 U7556 ( .IN(n3496), .QN(n1544) );
  AO222X1 U7557 ( .IN1(n4027), .IN2(n1730), .IN3(n4028), .IN4(g3227), .IN5(
        g3207), .IN6(n6114), .Q(g30401) );
  OA21X1 U7558 ( .IN1(n4017), .IN2(n3501), .IN3(n6372), .Q(n4028) );
  AO222X1 U7559 ( .IN1(n3931), .IN2(n6040), .IN3(n3932), .IN4(g5196), .IN5(
        g5188), .IN6(n6110), .Q(g30460) );
  NOR2X0 U7560 ( .IN1(n3931), .IN2(n6076), .QN(n3932) );
  ISOLANDX1 U7561 ( .D(n3926), .ISO(n3907), .Q(n3931) );
  AO222X1 U7562 ( .IN1(n3819), .IN2(n1511), .IN3(n3821), .IN4(g6271), .IN5(
        g6247), .IN6(n6089), .Q(g30529) );
  OA21X1 U7563 ( .IN1(n3802), .IN2(n3417), .IN3(n6396), .Q(n3821) );
  AO222X1 U7564 ( .IN1(n3995), .IN2(n1680), .IN3(n3996), .IN4(g3578), .IN5(
        g3558), .IN6(n6113), .Q(g30422) );
  OA21X1 U7565 ( .IN1(n3986), .IN2(n3492), .IN3(n6376), .Q(n3996) );
  AO222X1 U7566 ( .IN1(n3886), .IN2(n1969), .IN3(n3890), .IN4(g5571), .IN5(
        g5543), .IN6(n6094), .Q(g30485) );
  OA21X1 U7567 ( .IN1(n3874), .IN2(n3437), .IN3(n6387), .Q(n3890) );
  AO222X1 U7568 ( .IN1(n3984), .IN2(n1682), .IN3(n3988), .IN4(test_so43), 
        .IN5(g3586), .IN6(n6112), .Q(g30428) );
  OA21X1 U7569 ( .IN1(n3980), .IN2(n3489), .IN3(n6378), .Q(n3988) );
  AO222X1 U7570 ( .IN1(n3774), .IN2(n2225), .IN3(n3779), .IN4(g6641), .IN5(
        g6625), .IN6(n6103), .Q(g30556) );
  OA21X1 U7571 ( .IN1(n3404), .IN2(n3773), .IN3(n6402), .Q(n3779) );
  AO222X1 U7572 ( .IN1(n3793), .IN2(n6046), .IN3(n3794), .IN4(g6593), .IN5(
        g6597), .IN6(n6104), .Q(g30546) );
  NOR2X0 U7573 ( .IN1(n3793), .IN2(n6071), .QN(n3794) );
  ISOLANDX1 U7574 ( .D(n3792), .ISO(n3768), .Q(n3793) );
  AO222X1 U7575 ( .IN1(n3924), .IN2(n6040), .IN3(n3925), .IN4(g5216), .IN5(
        g5220), .IN6(n6096), .Q(g30463) );
  NOR2X0 U7576 ( .IN1(n3924), .IN2(n6076), .QN(n3925) );
  ISOLANDX1 U7577 ( .D(n3926), .ISO(n3910), .Q(n3924) );
  AO222X1 U7578 ( .IN1(n3948), .IN2(n6038), .IN3(n3949), .IN4(g3897), .IN5(
        test_so65), .IN6(n6111), .Q(g30452) );
  NOR2X0 U7579 ( .IN1(n3948), .IN2(n6076), .QN(n3949) );
  NOR2X0 U7580 ( .IN1(n3950), .IN2(n5648), .QN(n3948) );
  AO222X1 U7581 ( .IN1(n3785), .IN2(n2224), .IN3(n3786), .IN4(g6621), .IN5(
        g6601), .IN6(n6103), .Q(g30551) );
  OA21X1 U7582 ( .IN1(n3776), .IN2(n3407), .IN3(n6400), .Q(n3786) );
  AO222X1 U7583 ( .IN1(n3831), .IN2(n6044), .IN3(n3832), .IN4(g6235), .IN5(
        g6227), .IN6(n6089), .Q(g30523) );
  NOR2X0 U7584 ( .IN1(n3831), .IN2(n6072), .QN(n3832) );
  ISOLANDX1 U7585 ( .D(n3826), .ISO(n3807), .Q(n3831) );
  AO222X1 U7586 ( .IN1(n3951), .IN2(n1905), .IN3(n3954), .IN4(g3957), .IN5(
        g3941), .IN6(n6111), .Q(g30450) );
  OA21X1 U7587 ( .IN1(n3945), .IN2(n3479), .IN3(n6382), .Q(n3954) );
  AO222X1 U7588 ( .IN1(n3839), .IN2(n6043), .IN3(n3840), .IN4(g5897), .IN5(
        g5949), .IN6(n6090), .Q(g30518) );
  NOR2X0 U7589 ( .IN1(n3839), .IN2(n6072), .QN(n3840) );
  NOR2X0 U7590 ( .IN1(n3841), .IN2(n5649), .QN(n3839) );
  AO222X1 U7591 ( .IN1(n3908), .IN2(n1581), .IN3(n3909), .IN4(g5268), .IN5(
        g5252), .IN6(n6095), .Q(g30475) );
  OA21X1 U7592 ( .IN1(n3910), .IN2(n3444), .IN3(n6387), .Q(n3909) );
  AO222X1 U7593 ( .IN1(n3829), .IN2(n6043), .IN3(n3830), .IN4(g6239), .IN5(
        g6243), .IN6(n6089), .Q(g30524) );
  NOR2X0 U7594 ( .IN1(n3829), .IN2(n6072), .QN(n3830) );
  ISOLANDX1 U7595 ( .D(n3826), .ISO(n3804), .Q(n3829) );
  AO222X1 U7596 ( .IN1(n3819), .IN2(n1514), .IN3(n3820), .IN4(g6275), .IN5(
        g6255), .IN6(n6090), .Q(g30530) );
  OA21X1 U7597 ( .IN1(n3810), .IN2(n3417), .IN3(n6396), .Q(n3820) );
  AO222X1 U7598 ( .IN1(n3962), .IN2(n1904), .IN3(n3966), .IN4(g3917), .IN5(
        test_so24), .IN6(n6112), .Q(g30440) );
  OA21X1 U7599 ( .IN1(n3950), .IN2(n3482), .IN3(n6379), .Q(n3966) );
  AO222X1 U7600 ( .IN1(n3886), .IN2(n1970), .IN3(n3889), .IN4(g5575), .IN5(
        g5547), .IN6(n6094), .Q(g30486) );
  OA21X1 U7601 ( .IN1(n3871), .IN2(n3437), .IN3(n6387), .Q(n3889) );
  AO222X1 U7602 ( .IN1(n3842), .IN2(n1818), .IN3(n3845), .IN4(g5957), .IN5(
        g5941), .IN6(n6090), .Q(g30516) );
  OA21X1 U7603 ( .IN1(n3836), .IN2(n3424), .IN3(n6395), .Q(n3845) );
  AO222X1 U7604 ( .IN1(n3774), .IN2(n2226), .IN3(n3778), .IN4(g6645), .IN5(
        g6629), .IN6(n6103), .Q(g30557) );
  OA21X1 U7605 ( .IN1(n3770), .IN2(n3404), .IN3(n6402), .Q(n3778) );
  AO222X1 U7606 ( .IN1(n3951), .IN2(n1908), .IN3(n3952), .IN4(g3961), .IN5(
        g3945), .IN6(n6111), .Q(g30451) );
  OA21X1 U7607 ( .IN1(n3953), .IN2(n3479), .IN3(n6382), .Q(n3952) );
  AO222X1 U7608 ( .IN1(n3853), .IN2(n1817), .IN3(n3857), .IN4(test_so28), 
        .IN5(g5889), .IN6(n6091), .Q(g30506) );
  OA21X1 U7609 ( .IN1(n3841), .IN2(n3427), .IN3(n6391), .Q(n3857) );
  AO222X1 U7610 ( .IN1(n3886), .IN2(n1967), .IN3(n3888), .IN4(g5579), .IN5(
        g5555), .IN6(n6094), .Q(g30487) );
  OA21X1 U7611 ( .IN1(n3869), .IN2(n3437), .IN3(n6388), .Q(n3888) );
  AO222X1 U7612 ( .IN1(n3927), .IN2(n6040), .IN3(n3928), .IN4(g5208), .IN5(
        g5212), .IN6(n6096), .Q(g30462) );
  NOR2X0 U7613 ( .IN1(n3927), .IN2(n6063), .QN(n3928) );
  ISOLANDX1 U7614 ( .D(n3926), .ISO(n3902), .Q(n3927) );
  AO222X1 U7615 ( .IN1(n3774), .IN2(n2222), .IN3(n3777), .IN4(g6649), .IN5(
        g6633), .IN6(n6103), .Q(g30558) );
  OA21X1 U7616 ( .IN1(n3768), .IN2(n3404), .IN3(n6403), .Q(n3777) );
  AO222X1 U7617 ( .IN1(n3780), .IN2(n2226), .IN3(n3783), .IN4(g6629), .IN5(
        g6613), .IN6(n6103), .Q(g30553) );
  OA21X1 U7618 ( .IN1(n3770), .IN2(n3406), .IN3(n6401), .Q(n3783) );
  AO222X1 U7619 ( .IN1(n3974), .IN2(n6037), .IN3(n3975), .IN4(test_so24), 
        .IN5(g3881), .IN6(n6112), .Q(g30436) );
  NOR2X0 U7620 ( .IN1(n3974), .IN2(n6075), .QN(n3975) );
  ISOLANDX1 U7621 ( .D(n3969), .ISO(n3950), .Q(n3974) );
  AO222X1 U7622 ( .IN1(n3805), .IN2(n6044), .IN3(n3806), .IN4(g6243), .IN5(
        g6295), .IN6(n6105), .Q(g30539) );
  NOR2X0 U7623 ( .IN1(n3805), .IN2(n6072), .QN(n3806) );
  NOR2X0 U7624 ( .IN1(n3807), .IN2(n5651), .QN(n3805) );
  AO222X1 U7625 ( .IN1(n3842), .IN2(n1821), .IN3(n3843), .IN4(g5961), .IN5(
        g5945), .IN6(n6090), .Q(g30517) );
  OA21X1 U7626 ( .IN1(n3844), .IN2(n3424), .IN3(n6395), .Q(n3843) );
  AO222X1 U7627 ( .IN1(n3898), .IN2(n6041), .IN3(n3899), .IN4(g5543), .IN5(
        g5535), .IN6(n6094), .Q(g30481) );
  NOR2X0 U7628 ( .IN1(n3898), .IN2(n6075), .QN(n3899) );
  ISOLANDX1 U7629 ( .D(n3893), .ISO(n3874), .Q(n3898) );
  AO222X1 U7630 ( .IN1(n3995), .IN2(n1678), .IN3(n3997), .IN4(g3574), .IN5(
        g3550), .IN6(n6113), .Q(g30421) );
  OA21X1 U7631 ( .IN1(n3978), .IN2(n3492), .IN3(n6375), .Q(n3997) );
  AO222X1 U7632 ( .IN1(n3410), .IN2(n6045), .IN3(n3803), .IN4(g6251), .IN5(
        g6299), .IN6(n6105), .Q(g30540) );
  NOR2X0 U7633 ( .IN1(n3410), .IN2(n6072), .QN(n3803) );
  AO222X1 U7634 ( .IN1(n3970), .IN2(n6039), .IN3(n3971), .IN4(g3901), .IN5(
        g3905), .IN6(n6112), .Q(g30438) );
  NOR2X0 U7635 ( .IN1(n3970), .IN2(n6075), .QN(n3971) );
  ISOLANDX1 U7636 ( .D(n3969), .ISO(n3945), .Q(n3970) );
  AO222X1 U7637 ( .IN1(n4000), .IN2(n6036), .IN3(n4001), .IN4(g3558), .IN5(
        g3562), .IN6(n6113), .Q(g30418) );
  NOR2X0 U7638 ( .IN1(n4000), .IN2(n6074), .QN(n4001) );
  ISOLANDX1 U7639 ( .D(n4002), .ISO(n3986), .Q(n4000) );
  AO222X1 U7640 ( .IN1(n3872), .IN2(n6042), .IN3(n3873), .IN4(g5551), .IN5(
        g5603), .IN6(n6092), .Q(g30497) );
  NOR2X0 U7641 ( .IN1(n3872), .IN2(n6074), .QN(n3873) );
  NOR2X0 U7642 ( .IN1(n3874), .IN2(n5647), .QN(n3872) );
  AO222X1 U7643 ( .IN1(n3808), .IN2(n1514), .IN3(n3809), .IN4(g6307), .IN5(
        g6291), .IN6(n6105), .Q(g30538) );
  OA21X1 U7644 ( .IN1(n3810), .IN2(n3414), .IN3(n6399), .Q(n3809) );
  AO222X1 U7645 ( .IN1(n3780), .IN2(n2224), .IN3(n3781), .IN4(g6637), .IN5(
        g6621), .IN6(n6103), .Q(g30555) );
  OA21X1 U7646 ( .IN1(n3776), .IN2(n3406), .IN3(n6401), .Q(n3781) );
  AO222X1 U7647 ( .IN1(n3865), .IN2(n6042), .IN3(n3866), .IN4(g5889), .IN5(
        test_so36), .IN6(n6092), .Q(g30502) );
  NOR2X0 U7648 ( .IN1(n3865), .IN2(n6073), .QN(n3866) );
  ISOLANDX1 U7649 ( .D(n3860), .ISO(n3841), .Q(n3865) );
  AO222X1 U7650 ( .IN1(n3861), .IN2(n6043), .IN3(n3862), .IN4(g5901), .IN5(
        g5905), .IN6(n6091), .Q(g30504) );
  NOR2X0 U7651 ( .IN1(n3861), .IN2(n6073), .QN(n3862) );
  ISOLANDX1 U7652 ( .D(n3860), .ISO(n3836), .Q(n3861) );
  AO222X1 U7653 ( .IN1(n3995), .IN2(n1681), .IN3(n3999), .IN4(g3566), .IN5(
        g3538), .IN6(n6113), .Q(g30419) );
  OA21X1 U7654 ( .IN1(n3983), .IN2(n3492), .IN3(n6375), .Q(n3999) );
  AO222X1 U7655 ( .IN1(n4022), .IN2(n1732), .IN3(n4025), .IN4(g3235), .IN5(
        g3219), .IN6(n6115), .Q(g30403) );
  OA21X1 U7656 ( .IN1(n4020), .IN2(n3502), .IN3(n6372), .Q(n4025) );
  AO222X1 U7657 ( .IN1(n3875), .IN2(n1967), .IN3(n3878), .IN4(g5611), .IN5(
        g5595), .IN6(n6093), .Q(g30495) );
  OA21X1 U7658 ( .IN1(n3869), .IN2(n3434), .IN3(n6390), .Q(n3878) );
  AO222X1 U7659 ( .IN1(n3908), .IN2(n1578), .IN3(n3911), .IN4(g5264), .IN5(
        g5248), .IN6(n6095), .Q(g30474) );
  OA21X1 U7660 ( .IN1(n3902), .IN2(n3444), .IN3(n6386), .Q(n3911) );
  AO222X1 U7661 ( .IN1(n3819), .IN2(n1509), .IN3(n3822), .IN4(g6267), .IN5(
        g6239), .IN6(n6090), .Q(g30528) );
  OA21X1 U7662 ( .IN1(n3804), .IN2(n3417), .IN3(n6396), .Q(n3822) );
  AO222X1 U7663 ( .IN1(n3867), .IN2(n6042), .IN3(n3868), .IN4(g5567), .IN5(
        g5611), .IN6(n6092), .Q(g30499) );
  NOR2X0 U7664 ( .IN1(n3867), .IN2(n6073), .QN(n3868) );
  NOR2X0 U7665 ( .IN1(n3869), .IN2(n5647), .QN(n3867) );
  AO222X1 U7666 ( .IN1(n3824), .IN2(n6044), .IN3(n3825), .IN4(g6255), .IN5(
        g6259), .IN6(n6089), .Q(g30526) );
  NOR2X0 U7667 ( .IN1(n3824), .IN2(n6072), .QN(n3825) );
  ISOLANDX1 U7668 ( .D(n3826), .ISO(n3810), .Q(n3824) );
  AO222X1 U7669 ( .IN1(n3475), .IN2(n6039), .IN3(n3946), .IN4(g3905), .IN5(
        g3953), .IN6(n6111), .Q(g30453) );
  NOR2X0 U7670 ( .IN1(n3475), .IN2(n6076), .QN(n3946) );
  AO222X1 U7671 ( .IN1(n3894), .IN2(n6041), .IN3(n3895), .IN4(g5555), .IN5(
        test_so6), .IN6(n6105), .Q(g30483) );
  NOR2X0 U7672 ( .IN1(n3894), .IN2(n6074), .QN(n3895) );
  ISOLANDX1 U7673 ( .D(n3893), .ISO(n3869), .Q(n3894) );
  AO222X1 U7674 ( .IN1(n3995), .IN2(n1682), .IN3(n3998), .IN4(g3570), .IN5(
        g3542), .IN6(n6113), .Q(g30420) );
  OA21X1 U7675 ( .IN1(n3980), .IN2(n3492), .IN3(n6375), .Q(n3998) );
  AO222X1 U7676 ( .IN1(n3990), .IN2(n1682), .IN3(n3993), .IN4(g3586), .IN5(
        g3570), .IN6(n6113), .Q(g30424) );
  OA21X1 U7677 ( .IN1(n3980), .IN2(n3491), .IN3(n6376), .Q(n3993) );
  AO222X1 U7678 ( .IN1(n3984), .IN2(n1678), .IN3(n3987), .IN4(g3606), .IN5(
        g3590), .IN6(n6112), .Q(g30429) );
  OA21X1 U7679 ( .IN1(n3978), .IN2(n3489), .IN3(n6378), .Q(n3987) );
  AO222X1 U7680 ( .IN1(n3905), .IN2(n6040), .IN3(n3906), .IN4(g5204), .IN5(
        g5256), .IN6(n6095), .Q(g30476) );
  NOR2X0 U7681 ( .IN1(n3905), .IN2(n6076), .QN(n3906) );
  NOR2X0 U7682 ( .IN1(n3907), .IN2(n5650), .QN(n3905) );
  AO222X1 U7683 ( .IN1(n3420), .IN2(n6039), .IN3(n3837), .IN4(g5905), .IN5(
        g5953), .IN6(n6090), .Q(g30519) );
  NOR2X0 U7684 ( .IN1(n3420), .IN2(n6072), .QN(n3837) );
  AO222X1 U7685 ( .IN1(n3800), .IN2(n6045), .IN3(n3801), .IN4(g6259), .IN5(
        g6303), .IN6(n6105), .Q(g30541) );
  NOR2X0 U7686 ( .IN1(n3800), .IN2(n6072), .QN(n3801) );
  NOR2X0 U7687 ( .IN1(n3802), .IN2(n5651), .QN(n3800) );
  AO222X1 U7688 ( .IN1(n3967), .IN2(n6038), .IN3(n3968), .IN4(g3909), .IN5(
        g3913), .IN6(n6112), .Q(g30439) );
  NOR2X0 U7689 ( .IN1(n3967), .IN2(n6075), .QN(n3968) );
  ISOLANDX1 U7690 ( .D(n3969), .ISO(n3953), .Q(n3967) );
  AO222X1 U7691 ( .IN1(n3430), .IN2(n6042), .IN3(n3870), .IN4(test_so6), .IN5(
        g5607), .IN6(n6092), .Q(g30498) );
  NOR2X0 U7692 ( .IN1(n3430), .IN2(n6074), .QN(n3870) );
  AO222X1 U7693 ( .IN1(n3814), .IN2(n1514), .IN3(n3815), .IN4(g6291), .IN5(
        g6275), .IN6(n6089), .Q(g30534) );
  OA21X1 U7694 ( .IN1(n3810), .IN2(n3416), .IN3(n6397), .Q(n3815) );
  AO222X1 U7695 ( .IN1(n3984), .IN2(n1681), .IN3(n3989), .IN4(g3598), .IN5(
        g3582), .IN6(n6112), .Q(g30427) );
  OA21X1 U7696 ( .IN1(n3489), .IN2(n3983), .IN3(n6377), .Q(n3989) );
  AO222X1 U7697 ( .IN1(n3881), .IN2(n1970), .IN3(n3884), .IN4(test_so5), .IN5(
        g5575), .IN6(n6093), .Q(g30490) );
  OA21X1 U7698 ( .IN1(n3871), .IN2(n3436), .IN3(n6389), .Q(n3884) );
  AO222X1 U7699 ( .IN1(n3875), .IN2(n1968), .IN3(n3876), .IN4(g5615), .IN5(
        g5599), .IN6(n6093), .Q(g30496) );
  OA21X1 U7700 ( .IN1(n3877), .IN2(n3434), .IN3(n6391), .Q(n3876) );
  AO222X1 U7701 ( .IN1(n3875), .IN2(n1970), .IN3(n3879), .IN4(g5607), .IN5(
        test_so5), .IN6(n6093), .Q(g30494) );
  OA21X1 U7702 ( .IN1(n3871), .IN2(n3434), .IN3(n6390), .Q(n3879) );
  AO222X1 U7703 ( .IN1(n3485), .IN2(n6037), .IN3(n3979), .IN4(g3554), .IN5(
        test_so43), .IN6(n6112), .Q(g30432) );
  NOR2X0 U7704 ( .IN1(n3485), .IN2(n6075), .QN(n3979) );
  AO222X1 U7705 ( .IN1(n3858), .IN2(n6043), .IN3(n3859), .IN4(g5909), .IN5(
        g5913), .IN6(n6091), .Q(g30505) );
  NOR2X0 U7706 ( .IN1(n3858), .IN2(n6073), .QN(n3859) );
  ISOLANDX1 U7707 ( .D(n3860), .ISO(n3844), .Q(n3858) );
  AO222X1 U7708 ( .IN1(n3919), .IN2(n1578), .IN3(n3921), .IN4(g5232), .IN5(
        g5208), .IN6(n6096), .Q(g30466) );
  OA21X1 U7709 ( .IN1(n3902), .IN2(n3447), .IN3(n6384), .Q(n3921) );
  AO222X1 U7710 ( .IN1(n4005), .IN2(n6038), .IN3(n4006), .IN4(g3542), .IN5(
        g3546), .IN6(n6113), .Q(g30416) );
  NOR2X0 U7711 ( .IN1(n4005), .IN2(n6074), .QN(n4006) );
  ISOLANDX1 U7712 ( .D(n4002), .ISO(n3980), .Q(n4005) );
  AO222X1 U7713 ( .IN1(n4022), .IN2(n1730), .IN3(n4023), .IN4(g3243), .IN5(
        g3227), .IN6(n6114), .Q(g30405) );
  OA21X1 U7714 ( .IN1(n4017), .IN2(n3502), .IN3(n6373), .Q(n4023) );
  AO222X1 U7715 ( .IN1(n3881), .IN2(n1967), .IN3(n3883), .IN4(g5595), .IN5(
        g5579), .IN6(n6093), .Q(g30491) );
  OA21X1 U7716 ( .IN1(n3869), .IN2(n3436), .IN3(n6389), .Q(n3883) );
  AO222X1 U7717 ( .IN1(n3914), .IN2(n1578), .IN3(n3916), .IN4(g5248), .IN5(
        g5232), .IN6(n6096), .Q(g30470) );
  OA21X1 U7718 ( .IN1(n3902), .IN2(n3446), .IN3(n6385), .Q(n3916) );
  AO222X1 U7719 ( .IN1(n3957), .IN2(n1905), .IN3(n3959), .IN4(g3941), .IN5(
        g3925), .IN6(n6111), .Q(g30446) );
  OA21X1 U7720 ( .IN1(n3945), .IN2(n3481), .IN3(n6381), .Q(n3959) );
  AO222X1 U7721 ( .IN1(n3780), .IN2(n2222), .IN3(n3782), .IN4(g6633), .IN5(
        g6617), .IN6(n6103), .Q(g30554) );
  OA21X1 U7722 ( .IN1(n3768), .IN2(n3406), .IN3(n6402), .Q(n3782) );
  AO222X1 U7723 ( .IN1(n3848), .IN2(n1818), .IN3(n3850), .IN4(g5941), .IN5(
        g5925), .IN6(n6090), .Q(g30512) );
  OA21X1 U7724 ( .IN1(n3836), .IN2(n3426), .IN3(n6393), .Q(n3850) );
  AO222X1 U7725 ( .IN1(n3990), .IN2(n1678), .IN3(n3992), .IN4(g3590), .IN5(
        g3574), .IN6(n6113), .Q(g30425) );
  OA21X1 U7726 ( .IN1(n3978), .IN2(n3491), .IN3(n6377), .Q(n3992) );
  AO222X1 U7727 ( .IN1(n3914), .IN2(n1577), .IN3(n3918), .IN4(g5240), .IN5(
        g5224), .IN6(n6096), .Q(g30468) );
  OA21X1 U7728 ( .IN1(n3446), .IN2(n3907), .IN3(n6384), .Q(n3918) );
  AO222X1 U7729 ( .IN1(n3990), .IN2(n1681), .IN3(n3994), .IN4(g3582), .IN5(
        g3566), .IN6(n6113), .Q(g30423) );
  OA21X1 U7730 ( .IN1(n3491), .IN2(n3983), .IN3(n6376), .Q(n3994) );
  AO222X1 U7731 ( .IN1(n3780), .IN2(n2225), .IN3(n3784), .IN4(g6625), .IN5(
        g6609), .IN6(n6103), .Q(g30552) );
  OA21X1 U7732 ( .IN1(n3406), .IN2(n3773), .IN3(n6401), .Q(n3784) );
  AO222X1 U7733 ( .IN1(n3814), .IN2(n1510), .IN3(n3818), .IN4(g6279), .IN5(
        g6263), .IN6(n6089), .Q(g30531) );
  OA21X1 U7734 ( .IN1(n3416), .IN2(n3807), .IN3(n6397), .Q(n3818) );
  AO222X1 U7735 ( .IN1(n4022), .IN2(n1731), .IN3(n4026), .IN4(g3231), .IN5(
        g3215), .IN6(n6115), .Q(g30402) );
  OA21X1 U7736 ( .IN1(n3502), .IN2(n4014), .IN3(n6394), .Q(n4026) );
  AO222X1 U7737 ( .IN1(n3957), .IN2(n1904), .IN3(n3961), .IN4(g3933), .IN5(
        g3917), .IN6(n6111), .Q(g30444) );
  OA21X1 U7738 ( .IN1(n3481), .IN2(n3950), .IN3(n6380), .Q(n3961) );
  AO222X1 U7739 ( .IN1(n3848), .IN2(n1817), .IN3(n3852), .IN4(g5933), .IN5(
        test_so28), .IN6(n6091), .Q(g30510) );
  OA21X1 U7740 ( .IN1(n3426), .IN2(n3841), .IN3(n6392), .Q(n3852) );
  AO222X1 U7741 ( .IN1(n4022), .IN2(n1729), .IN3(n4024), .IN4(g3239), .IN5(
        g3223), .IN6(n6114), .Q(g30404) );
  OA21X1 U7742 ( .IN1(n3502), .IN2(n3495), .IN3(n6373), .Q(n4024) );
  AO222X1 U7743 ( .IN1(n3814), .IN2(n1511), .IN3(n3816), .IN4(g6287), .IN5(
        g6271), .IN6(n6089), .Q(g30533) );
  OA21X1 U7744 ( .IN1(n3802), .IN2(n3416), .IN3(n6398), .Q(n3816) );
  AO222X1 U7745 ( .IN1(n3881), .IN2(n1969), .IN3(n3885), .IN4(g5587), .IN5(
        g5571), .IN6(n6093), .Q(g30489) );
  OA21X1 U7746 ( .IN1(n3436), .IN2(n3874), .IN3(n6388), .Q(n3885) );
  AO222X1 U7747 ( .IN1(n4863), .IN2(n1648), .IN3(n4866), .IN4(g4375), .IN5(
        g4411), .IN6(n6109), .Q(g26945) );
  AO222X1 U7748 ( .IN1(n2419), .IN2(n5291), .IN3(n2424), .IN4(n2404), .IN5(
        g790), .IN6(n6096), .Q(g34850) );
  NOR2X0 U7749 ( .IN1(n2419), .IN2(n5291), .QN(n2424) );
  AO222X1 U7750 ( .IN1(n2405), .IN2(n5479), .IN3(n2418), .IN4(n2404), .IN5(
        g794), .IN6(n6096), .Q(g34881) );
  NOR2X0 U7751 ( .IN1(n2405), .IN2(n5479), .QN(n2418) );
  AO222X1 U7752 ( .IN1(n6036), .IN2(g32975), .IN3(g5272), .IN4(n1434), .IN5(
        g5268), .IN6(n6095), .Q(g30479) );
  AO222X1 U7753 ( .IN1(n2404), .IN2(g554), .IN3(n2405), .IN4(g807), .IN5(g807), 
        .IN6(n6097), .Q(g34911) );
  NOR2X0 U7754 ( .IN1(g34975), .IN2(n6076), .QN(n2493) );
  AO222X1 U7755 ( .IN1(n6035), .IN2(n1546), .IN3(g3263), .IN4(n1440), .IN5(
        test_so84), .IN6(n6113), .Q(g30413) );
  AO222X1 U7756 ( .IN1(n6036), .IN2(n1755), .IN3(g5619), .IN4(n1433), .IN5(
        g5615), .IN6(n6092), .Q(g30500) );
  AO222X1 U7757 ( .IN1(n6036), .IN2(n1679), .IN3(g3614), .IN4(n1439), .IN5(
        g3610), .IN6(n6112), .Q(g30434) );
  AO222X1 U7758 ( .IN1(n6035), .IN2(n2223), .IN3(g6657), .IN4(n1430), .IN5(
        g6653), .IN6(n6102), .Q(g30563) );
  AO222X1 U7759 ( .IN1(n6035), .IN2(n1513), .IN3(g6311), .IN4(n1431), .IN5(
        g6307), .IN6(n6104), .Q(g30542) );
  AO222X1 U7760 ( .IN1(n6035), .IN2(n1907), .IN3(g3965), .IN4(n1438), .IN5(
        g3961), .IN6(n6110), .Q(g30455) );
  AO222X1 U7761 ( .IN1(n6035), .IN2(n1820), .IN3(test_so13), .IN4(n1432), 
        .IN5(g5961), .IN6(n6090), .Q(g30521) );
  OA21X1 U7762 ( .IN1(g6191), .IN2(g6177), .IN3(n6372), .Q(n4848) );
  OR2X1 U7763 ( .IN1(n5121), .IN2(g370), .Q(n4824) );
  AO22X1 U7764 ( .IN1(n1648), .IN2(n4864), .IN3(g4375), .IN4(n4865), .Q(g26946) );
  AO22X1 U7765 ( .IN1(n6134), .IN2(g550), .IN3(g21292), .IN4(n6289), .Q(g34598) );
  AO221X1 U7766 ( .IN1(n3628), .IN2(g1783), .IN3(g1798), .IN4(n6085), .IN5(
        n3629), .Q(g32993) );
  AO21X1 U7767 ( .IN1(n1397), .IN2(g1792), .IN3(n3630), .Q(n3629) );
  AO221X1 U7768 ( .IN1(n3593), .IN2(g2051), .IN3(g2066), .IN4(n6085), .IN5(
        n3594), .Q(g33001) );
  AO21X1 U7769 ( .IN1(n1395), .IN2(g2060), .IN3(n3595), .Q(n3594) );
  AO221X1 U7770 ( .IN1(n3574), .IN2(g2208), .IN3(g2223), .IN4(n6086), .IN5(
        n3575), .Q(g33005) );
  AO21X1 U7771 ( .IN1(n1394), .IN2(g2217), .IN3(n3576), .Q(n3575) );
  AO221X1 U7772 ( .IN1(n3555), .IN2(test_so21), .IN3(g2357), .IN4(n6086), 
        .IN5(n3556), .Q(g33009) );
  AO21X1 U7773 ( .IN1(n1393), .IN2(g2351), .IN3(n3557), .Q(n3556) );
  AO221X1 U7774 ( .IN1(n3517), .IN2(g2610), .IN3(test_so40), .IN4(n6087), 
        .IN5(n3518), .Q(g33017) );
  AO21X1 U7775 ( .IN1(n1391), .IN2(g2619), .IN3(n3519), .Q(n3518) );
  AO221X1 U7776 ( .IN1(n3536), .IN2(g2476), .IN3(g2491), .IN4(n6086), .IN5(
        n3537), .Q(g33013) );
  AO21X1 U7777 ( .IN1(n1392), .IN2(g2485), .IN3(n3538), .Q(n3537) );
  AO221X1 U7778 ( .IN1(n3611), .IN2(g1917), .IN3(g1932), .IN4(n6086), .IN5(
        n3612), .Q(g32997) );
  AO21X1 U7779 ( .IN1(n1396), .IN2(g1926), .IN3(n3613), .Q(n3612) );
  AO221X1 U7780 ( .IN1(n3646), .IN2(test_so94), .IN3(g1664), .IN4(n6086), 
        .IN5(n3647), .Q(g32989) );
  AO21X1 U7781 ( .IN1(n1398), .IN2(g1657), .IN3(n3648), .Q(n3647) );
  OR2X1 U7782 ( .IN1(n3648), .IN2(n5973), .Q(n3650) );
  AND3X1 U7783 ( .IN1(n3652), .IN2(n5525), .IN3(n3646), .Q(n5973) );
  OR2X1 U7784 ( .IN1(n3630), .IN2(n5974), .Q(n3632) );
  AND3X1 U7785 ( .IN1(n3634), .IN2(n5359), .IN3(n3628), .Q(n5974) );
  OA21X1 U7786 ( .IN1(test_so83), .IN2(g5831), .IN3(n6360), .Q(n4846) );
  NAND2X0 U7787 ( .IN1(g5817), .IN2(n6158), .QN(n3760) );
  NAND2X0 U7788 ( .IN1(g6163), .IN2(n6172), .QN(n3761) );
  AO22X1 U7789 ( .IN1(n6274), .IN2(g4411), .IN3(n4873), .IN4(g4401), .Q(g26949) );
  AO21X1 U7790 ( .IN1(g4392), .IN2(n1648), .IN3(n6137), .Q(n4873) );
  AO21X1 U7791 ( .IN1(g947), .IN2(n6122), .IN3(n2504), .Q(g34726) );
  ISOLANDX1 U7792 ( .D(g952), .ISO(n6145), .Q(n2505) );
  AO21X1 U7793 ( .IN1(g1291), .IN2(n6121), .IN3(n2498), .Q(g34729) );
  ISOLANDX1 U7794 ( .D(g1296), .ISO(n6144), .Q(n2499) );
  AO21X1 U7795 ( .IN1(g538), .IN2(n6122), .IN3(n2512), .Q(g34722) );
  AO21X1 U7796 ( .IN1(g2856), .IN2(n6120), .IN3(n2472), .Q(g34794) );
  AO21X1 U7797 ( .IN1(g2917), .IN2(n6120), .IN3(n2450), .Q(g34803) );
  OR2X1 U7798 ( .IN1(g2927), .IN2(g2932), .Q(n2451) );
  XNOR2X1 U7799 ( .IN1(g4332), .IN2(n6016), .Q(n3060) );
  AO21X1 U7800 ( .IN1(g939), .IN2(n6122), .IN3(n2500), .Q(g34728) );
  NOR2X0 U7801 ( .IN1(n5409), .IN2(n6076), .QN(n2502) );
  AO21X1 U7802 ( .IN1(g1283), .IN2(n6122), .IN3(n2494), .Q(g34731) );
  NOR2X0 U7803 ( .IN1(n5623), .IN2(n6077), .QN(n2496) );
  AO22X1 U7804 ( .IN1(g2955), .IN2(n6123), .IN3(n2429), .IN4(n6276), .Q(g34808) );
  OR4X1 U7805 ( .IN1(n5926), .IN2(n2432), .IN3(n2433), .IN4(g2965), .Q(n2429)
         );
  NAND2X0 U7806 ( .IN1(g5471), .IN2(n6160), .QN(n3758) );
  OR4X1 U7807 ( .IN1(n2393), .IN2(g24161), .IN3(g24162), .IN4(g24163), .Q(
        n2397) );
  NBUFFX2 U7808 ( .IN(g72), .Q(g24166) );
  NOR2X0 U7809 ( .IN1(n2549), .IN2(n6078), .QN(g34602) );
  NBUFFX2 U7810 ( .IN(g73), .Q(n6016) );
  AOI21X1 U7811 ( .IN1(g12184), .IN2(n5482), .IN3(n4205), .QN(n4199) );
  NAND2X0 U7812 ( .IN1(n2394), .IN2(n2395), .QN(g34980) );
  NAND2X0 U7813 ( .IN1(test_so14), .IN2(n6079), .QN(n2394) );
  OA221X1 U7814 ( .IN1(n6026), .IN2(n5975), .IN3(n6026), .IN4(n5976), .IN5(
        n3333), .Q(n3387) );
  AOI221X1 U7815 ( .IN1(g2890), .IN2(n1800), .IN3(g24173), .IN4(n1801), .IN5(
        n3393), .QN(n5975) );
  AOI221X1 U7816 ( .IN1(test_so60), .IN2(n1788), .IN3(g199), .IN4(n1790), 
        .IN5(n3390), .QN(n5976) );
  NOR2X0 U7817 ( .IN1(g2724), .IN2(g2729), .QN(n4062) );
  NAND2X0 U7818 ( .IN1(g2719), .IN2(g2715), .QN(n4052) );
  NAND4X0 U7819 ( .IN1(n2994), .IN2(n2995), .IN3(n2996), .IN4(n2997), .QN(
        g34781) );
  OA22X1 U7820 ( .IN1(n5596), .IN2(n3002), .IN3(n3003), .IN4(n3004), .Q(n2996)
         );
  NAND3X0 U7821 ( .IN1(n1467), .IN2(n5510), .IN3(g1917), .QN(n2994) );
  NAND3X0 U7822 ( .IN1(n1468), .IN2(n5507), .IN3(g2051), .QN(n2995) );
  NAND2X0 U7823 ( .IN1(g12919), .IN2(n6173), .QN(n3269) );
  NAND2X0 U7824 ( .IN1(g12923), .IN2(n6156), .QN(n3261) );
  NAND2X0 U7825 ( .IN1(g2719), .IN2(n5299), .QN(n4051) );
  AO221X1 U7826 ( .IN1(n3197), .IN2(g2130), .IN3(g956), .IN4(n5286), .IN5(
        n2978), .Q(n2892) );
  NOR2X0 U7827 ( .IN1(n5275), .IN2(n5307), .QN(n3197) );
  AO221X1 U7828 ( .IN1(n3253), .IN2(g2130), .IN3(g1135), .IN4(n5286), .IN5(
        n2978), .Q(n2962) );
  NOR2X0 U7829 ( .IN1(g2145), .IN2(g2138), .QN(n3253) );
  AO221X1 U7830 ( .IN1(n3236), .IN2(g2130), .IN3(g1105), .IN4(n5286), .IN5(
        n2978), .Q(n2939) );
  NOR2X0 U7831 ( .IN1(g2138), .IN2(n5307), .QN(n3236) );
  AO221X1 U7832 ( .IN1(n3217), .IN2(g2130), .IN3(g1129), .IN4(n5286), .IN5(
        n2978), .Q(n2916) );
  NOR2X0 U7833 ( .IN1(g2145), .IN2(n5275), .QN(n3217) );
  NOR2X0 U7834 ( .IN1(test_so25), .IN2(g19), .QN(n3381) );
  NAND2X0 U7835 ( .IN1(g1783), .IN2(n5602), .QN(n3634) );
  NOR2X0 U7836 ( .IN1(n6239), .IN2(DFF_1381_n1), .QN(g21727) );
  AND2X1 U7837 ( .IN1(g1536), .IN2(n4836), .Q(n3177) );
  OA21X1 U7838 ( .IN1(g5152), .IN2(g5138), .IN3(n6364), .Q(n2471) );
  AND2X1 U7839 ( .IN1(g1193), .IN2(n4837), .Q(n3254) );
  NAND2X0 U7840 ( .IN1(n2972), .IN2(g1668), .QN(n2971) );
  NOR2X0 U7841 ( .IN1(n2587), .IN2(g4639), .QN(g34025) );
  OA21X1 U7842 ( .IN1(g3494), .IN2(g3480), .IN3(n6354), .Q(n4852) );
  NAND2X0 U7843 ( .IN1(n2775), .IN2(test_so81), .QN(n2733) );
  NAND2X0 U7844 ( .IN1(n2761), .IN2(test_so81), .QN(n2740) );
  NAND2X0 U7845 ( .IN1(test_so79), .IN2(n2827), .QN(n2832) );
  NAND2X0 U7846 ( .IN1(g2153), .IN2(n2873), .QN(n2878) );
  NAND2X0 U7847 ( .IN1(g2555), .IN2(n2803), .QN(n2808) );
  NAND2X0 U7848 ( .IN1(g1996), .IN2(n2896), .QN(n2901) );
  NAND2X0 U7849 ( .IN1(g2287), .IN2(n2850), .QN(n2855) );
  NAND2X0 U7850 ( .IN1(g1728), .IN2(n2943), .QN(n2948) );
  NAND2X0 U7851 ( .IN1(test_so8), .IN2(n2920), .QN(n2925) );
  NAND2X0 U7852 ( .IN1(g20049), .IN2(n1402), .QN(n3463) );
  NAND2X0 U7853 ( .IN1(g4169), .IN2(n6176), .QN(n5027) );
  OA21X1 U7854 ( .IN1(n2892), .IN2(g23683), .IN3(n2893), .Q(n2886) );
  OA21X1 U7855 ( .IN1(n2939), .IN2(g23683), .IN3(n2940), .Q(n2933) );
  AO221X1 U7856 ( .IN1(n3137), .IN2(g2689), .IN3(g1472), .IN4(n2549), .IN5(
        n1342), .Q(n2822) );
  NOR2X0 U7857 ( .IN1(g2704), .IN2(n5308), .QN(n3137) );
  AO221X1 U7858 ( .IN1(n3176), .IN2(g2689), .IN3(g1478), .IN4(n2549), .IN5(
        n1342), .Q(n2868) );
  NOR2X0 U7859 ( .IN1(g2704), .IN2(g2697), .QN(n3176) );
  AO221X1 U7860 ( .IN1(n3118), .IN2(g2689), .IN3(g1300), .IN4(n2549), .IN5(
        n1342), .Q(n2798) );
  NOR2X0 U7861 ( .IN1(n5308), .IN2(n5377), .QN(n3118) );
  AO221X1 U7862 ( .IN1(n3156), .IN2(g2689), .IN3(g1448), .IN4(n2549), .IN5(
        n1342), .Q(n2845) );
  NOR2X0 U7863 ( .IN1(g2697), .IN2(n5377), .QN(n3156) );
  OA21X1 U7864 ( .IN1(n2798), .IN2(g1585), .IN3(n2799), .Q(n2792) );
  OA21X1 U7865 ( .IN1(n2845), .IN2(g1585), .IN3(n2846), .Q(n2839) );
  NOR2X0 U7866 ( .IN1(n5349), .IN2(g2748), .QN(n3562) );
  AND3X1 U7867 ( .IN1(n2531), .IN2(n3381), .IN3(g9), .Q(n2546) );
  AND3X1 U7868 ( .IN1(n3396), .IN2(n5469), .IN3(g28), .Q(n2528) );
  NOR2X0 U7869 ( .IN1(n5516), .IN2(g2741), .QN(n3543) );
  NOR2X0 U7870 ( .IN1(n6081), .IN2(g1306), .QN(n2447) );
  NAND3X0 U7871 ( .IN1(n1855), .IN2(g1792), .IN3(g1760), .QN(n4139) );
  NAND3X0 U7872 ( .IN1(n1745), .IN2(g2351), .IN3(g2319), .QN(n4091) );
  AO22X1 U7873 ( .IN1(g1848), .IN2(n4141), .IN3(n1409), .IN4(g1854), .Q(g30356) );
  INVX0 U7874 ( .IN(n4141), .QN(n1409) );
  NAND2X0 U7875 ( .IN1(n6213), .IN2(n4139), .QN(n4141) );
  AO22X1 U7876 ( .IN1(g1982), .IN2(n4129), .IN3(n1408), .IN4(g1988), .Q(g30361) );
  INVX0 U7877 ( .IN(n4129), .QN(n1408) );
  NAND2X0 U7878 ( .IN1(n6208), .IN2(n4127), .QN(n4129) );
  AO22X1 U7879 ( .IN1(g2675), .IN2(n4069), .IN3(n1403), .IN4(g2681), .Q(g30386) );
  INVX0 U7880 ( .IN(n4069), .QN(n1403) );
  NAND2X0 U7881 ( .IN1(n6195), .IN2(n4067), .QN(n4069) );
  AO22X1 U7882 ( .IN1(g1714), .IN2(n4153), .IN3(n1410), .IN4(g1720), .Q(g30351) );
  INVX0 U7883 ( .IN(n4153), .QN(n1410) );
  NAND2X0 U7884 ( .IN1(n6233), .IN2(n4151), .QN(n4153) );
  AO22X1 U7885 ( .IN1(g2273), .IN2(n4105), .IN3(n1406), .IN4(g2279), .Q(g30371) );
  INVX0 U7886 ( .IN(n4105), .QN(n1406) );
  NAND2X0 U7887 ( .IN1(n6199), .IN2(n4103), .QN(n4105) );
  AO22X1 U7888 ( .IN1(g2116), .IN2(n4117), .IN3(n1407), .IN4(g2122), .Q(g30366) );
  INVX0 U7889 ( .IN(n4117), .QN(n1407) );
  NAND2X0 U7890 ( .IN1(n6196), .IN2(n4115), .QN(n4117) );
  NOR2X0 U7891 ( .IN1(n5977), .IN2(n5978), .QN(n3581) );
  XOR2X1 U7892 ( .IN1(g2759), .IN2(n6018), .Q(n5977) );
  XOR2X1 U7893 ( .IN1(g2763), .IN2(n6016), .Q(n5978) );
  AND4X1 U7894 ( .IN1(g31), .IN2(g28), .IN3(n3396), .IN4(n5468), .Q(n3392) );
  ISOLANDX1 U7895 ( .D(n2668), .ISO(g24174), .Q(n2760) );
  AND4X1 U7896 ( .IN1(g9), .IN2(g8), .IN3(n3395), .IN4(test_so85), .Q(n3382)
         );
  ISOLANDX1 U7897 ( .D(g6), .ISO(g31), .Q(n3395) );
  NOR2X0 U7898 ( .IN1(n5477), .IN2(g19), .QN(n3394) );
  NAND2X0 U7899 ( .IN1(g4572), .IN2(n1402), .QN(n3462) );
  NAND2X0 U7900 ( .IN1(g4578), .IN2(n1402), .QN(n3453) );
  AND3X1 U7901 ( .IN1(n3750), .IN2(n1605), .IN3(test_so73), .Q(n3687) );
  AND3X1 U7902 ( .IN1(test_so55), .IN2(n1516), .IN3(test_so51), .Q(n3279) );
  NOR2X0 U7903 ( .IN1(n3348), .IN2(n3349), .QN(n3347) );
  AO221X1 U7904 ( .IN1(test_so95), .IN2(n2546), .IN3(g2941), .IN4(n2459), 
        .IN5(n3350), .Q(n3348) );
  AO222X1 U7905 ( .IN1(g2898), .IN2(n1793), .IN3(g2936), .IN4(n6001), .IN5(
        g2988), .IN6(n1800), .Q(n3349) );
  AND4X1 U7906 ( .IN1(n3382), .IN2(g19), .IN3(g28), .IN4(n5477), .Q(n3350) );
  AO22X1 U7907 ( .IN1(g6167), .IN2(n4231), .IN3(n1413), .IN4(g6173), .Q(g29300) );
  INVX0 U7908 ( .IN(n4231), .QN(n1413) );
  NAND2X0 U7909 ( .IN1(n6219), .IN2(n1566), .QN(n4231) );
  AO22X1 U7910 ( .IN1(g3821), .IN2(n4337), .IN3(n1418), .IN4(g3827), .Q(g29271) );
  INVX0 U7911 ( .IN(n4337), .QN(n1418) );
  NAND2X0 U7912 ( .IN1(n6228), .IN2(n1502), .QN(n4337) );
  AO22X1 U7913 ( .IN1(test_so96), .IN2(n4276), .IN3(n1416), .IN4(g5134), .Q(
        g29282) );
  INVX0 U7914 ( .IN(n4276), .QN(n1416) );
  NAND2X0 U7915 ( .IN1(n6234), .IN2(n1559), .QN(n4276) );
  AO22X1 U7916 ( .IN1(g3119), .IN2(n4367), .IN3(n1420), .IN4(g3125), .Q(g29259) );
  INVX0 U7917 ( .IN(n4367), .QN(n1420) );
  NAND2X0 U7918 ( .IN1(n6229), .IN2(n1589), .QN(n4367) );
  AO22X1 U7919 ( .IN1(g5475), .IN2(n4261), .IN3(n1415), .IN4(g5481), .Q(g29288) );
  INVX0 U7920 ( .IN(n4261), .QN(n1415) );
  NAND2X0 U7921 ( .IN1(n6220), .IN2(n1561), .QN(n4261) );
  AO22X1 U7922 ( .IN1(g5821), .IN2(n4246), .IN3(n1414), .IN4(g5827), .Q(g29294) );
  INVX0 U7923 ( .IN(n4246), .QN(n1414) );
  NAND2X0 U7924 ( .IN1(n6230), .IN2(n1563), .QN(n4246) );
  AO22X1 U7925 ( .IN1(g6513), .IN2(n4216), .IN3(n1412), .IN4(g6519), .Q(g29306) );
  INVX0 U7926 ( .IN(n4216), .QN(n1412) );
  NAND2X0 U7927 ( .IN1(n6205), .IN2(n1674), .QN(n4216) );
  AO22X1 U7928 ( .IN1(g3470), .IN2(n4352), .IN3(n1419), .IN4(g3476), .Q(g29265) );
  INVX0 U7929 ( .IN(n4352), .QN(n1419) );
  NAND2X0 U7930 ( .IN1(n6238), .IN2(n1594), .QN(n4352) );
  AND3X1 U7931 ( .IN1(n4204), .IN2(n4205), .IN3(g691), .Q(n3750) );
  NAND2X0 U7932 ( .IN1(n1605), .IN2(n4206), .QN(n4204) );
  NAND3X0 U7933 ( .IN1(n5402), .IN2(n5306), .IN3(n5606), .QN(n4206) );
  AO222X1 U7934 ( .IN1(g2970), .IN2(n6001), .IN3(g2975), .IN4(n2459), .IN5(
        g2886), .IN6(n1793), .Q(n3379) );
  NAND2X0 U7935 ( .IN1(g4180), .IN2(n2884), .QN(n2814) );
  AO222X1 U7936 ( .IN1(n1445), .IN2(g17423), .IN3(n5206), .IN4(g10527), .IN5(
        g1589), .IN6(n6108), .Q(g24255) );
  NOR2X0 U7937 ( .IN1(g17423), .IN2(n6078), .QN(n5206) );
  AO222X1 U7938 ( .IN1(n1447), .IN2(g17400), .IN3(n5228), .IN4(g10500), .IN5(
        g1246), .IN6(n6108), .Q(g24239) );
  NOR2X0 U7939 ( .IN1(g17400), .IN2(n6078), .QN(n5228) );
  NAND3X0 U7940 ( .IN1(g504), .IN2(g518), .IN3(n3195), .QN(n3206) );
  NAND3X0 U7941 ( .IN1(g504), .IN2(n5287), .IN3(n3195), .QN(n3226) );
  NAND3X0 U7942 ( .IN1(g518), .IN2(n5519), .IN3(n3195), .QN(n3186) );
  AND3X1 U7943 ( .IN1(n3396), .IN2(n5324), .IN3(g31), .Q(n3391) );
  AND3X1 U7944 ( .IN1(g19), .IN2(n5477), .IN3(g9), .Q(n3397) );
  NAND3X0 U7945 ( .IN1(n2528), .IN2(n3381), .IN3(g9), .QN(n3338) );
  NAND3X0 U7946 ( .IN1(n4830), .IN2(n4205), .IN3(g691), .QN(n3748) );
  OAI22X1 U7947 ( .IN1(n4834), .IN2(g278), .IN3(n5627), .IN4(n4835), .QN(n4830) );
  NAND3X0 U7948 ( .IN1(n1481), .IN2(n5505), .IN3(g2070), .QN(n2716) );
  NAND3X0 U7949 ( .IN1(n1479), .IN2(n5503), .IN3(g1936), .QN(n2715) );
  NAND3X0 U7950 ( .IN1(g1783), .IN2(n5359), .IN3(n1855), .QN(n4147) );
  NAND3X0 U7951 ( .IN1(test_so21), .IN2(n5511), .IN3(n1745), .QN(n4099) );
  NAND3X0 U7952 ( .IN1(n3116), .IN2(n5287), .IN3(g504), .QN(n3146) );
  NAND3X0 U7953 ( .IN1(n1477), .IN2(n5504), .IN3(g1802), .QN(n2725) );
  XNOR2X1 U7954 ( .IN1(n4497), .IN2(g1105), .Q(n4495) );
  XNOR2X1 U7955 ( .IN1(n4473), .IN2(g1300), .Q(n4478) );
  XNOR2X1 U7956 ( .IN1(n4473), .IN2(g1448), .Q(n4471) );
  AND3X1 U7957 ( .IN1(n1483), .IN2(n5513), .IN3(g2361), .Q(n2721) );
  XNOR2X1 U7958 ( .IN1(n4497), .IN2(g1135), .Q(n4512) );
  XNOR2X1 U7959 ( .IN1(n4497), .IN2(g956), .Q(n4502) );
  XNOR2X1 U7960 ( .IN1(n4497), .IN2(g1129), .Q(n4507) );
  XNOR2X1 U7961 ( .IN1(n4473), .IN2(g1472), .Q(n4483) );
  XNOR2X1 U7962 ( .IN1(n4473), .IN2(g1478), .Q(n4488) );
  AND3X1 U7963 ( .IN1(n1482), .IN2(n5514), .IN3(g2227), .Q(n2722) );
  AND3X1 U7964 ( .IN1(g996), .IN2(n6352), .IN3(n6021), .Q(n5078) );
  AO22X1 U7965 ( .IN1(g25219), .IN2(n6126), .IN3(n5159), .IN4(n6284), .Q(
        g24338) );
  NOR2X0 U7966 ( .IN1(g5352), .IN2(n5158), .QN(n5159) );
  AO22X1 U7967 ( .IN1(g25219), .IN2(n6272), .IN3(g5062), .IN4(n6136), .Q(
        g25701) );
  AND4X1 U7968 ( .IN1(n2998), .IN2(n2999), .IN3(n3000), .IN4(n3001), .Q(n2997)
         );
  NAND3X0 U7969 ( .IN1(n1470), .IN2(n5511), .IN3(test_so21), .QN(n2999) );
  NAND3X0 U7970 ( .IN1(n1471), .IN2(n5509), .IN3(g2476), .QN(n3000) );
  NAND3X0 U7971 ( .IN1(n1472), .IN2(n5508), .IN3(g2610), .QN(n3001) );
  NAND2X0 U7972 ( .IN1(g4581), .IN2(n6159), .QN(n3456) );
  NOR2X0 U7973 ( .IN1(g4382), .IN2(n6066), .QN(n4866) );
  AO222X1 U7974 ( .IN1(n1429), .IN2(g20899), .IN3(n4956), .IN4(n4532), .IN5(
        g728), .IN6(n4957), .Q(g26896) );
  INVX0 U7975 ( .IN(n4957), .QN(n1429) );
  NAND2X0 U7976 ( .IN1(n6217), .IN2(n1538), .QN(n4957) );
  ISOLANDX1 U7977 ( .D(g661), .ISO(n6145), .Q(n4956) );
  AO221X1 U7978 ( .IN1(g2955), .IN2(n2459), .IN3(g2950), .IN4(n6001), .IN5(
        n3350), .Q(n3360) );
  OA22X1 U7979 ( .IN1(n2731), .IN2(n5348), .IN3(g4358), .IN4(n2732), .Q(n2428)
         );
  OA221X1 U7980 ( .IN1(n2733), .IN2(n2734), .IN3(n2735), .IN4(n2736), .IN5(
        n2737), .Q(n2732) );
  OA221X1 U7981 ( .IN1(n2733), .IN2(n2742), .IN3(n2735), .IN4(n2743), .IN5(
        n2744), .Q(n2731) );
  OA22X1 U7982 ( .IN1(n2738), .IN2(n2739), .IN3(n2740), .IN4(n2741), .Q(n2737)
         );
  OA221X1 U7983 ( .IN1(g2994), .IN2(n3337), .IN3(n3338), .IN4(n5489), .IN5(
        n3339), .Q(n3334) );
  AOI222X1 U7984 ( .IN1(n6001), .IN2(g2922), .IN3(n2546), .IN4(g2860), .IN5(
        n2459), .IN6(g2927), .QN(n3339) );
  AO22X1 U7985 ( .IN1(g29218), .IN2(n6126), .IN3(n5163), .IN4(n5164), .Q(
        g24335) );
  NOR2X0 U7986 ( .IN1(g4340), .IN2(n5382), .QN(n5163) );
  OA221X1 U7987 ( .IN1(n3311), .IN2(n5491), .IN3(n3312), .IN4(n5330), .IN5(
        n3313), .Q(n3310) );
  OA22X1 U7988 ( .IN1(n3314), .IN2(n5476), .IN3(n3315), .IN4(n5338), .Q(n3313)
         );
  OA21X1 U7989 ( .IN1(g5499), .IN2(g5485), .IN3(n6353), .Q(n4843) );
  AO222X1 U7990 ( .IN1(g599), .IN2(n1794), .IN3(g562), .IN4(n1795), .IN5(g781), 
        .IN6(n1791), .Q(n3390) );
  AOI221X1 U7991 ( .IN1(n1800), .IN2(g2999), .IN3(n1793), .IN4(g2856), .IN5(
        n3328), .QN(n3326) );
  AO222X1 U7992 ( .IN1(n6001), .IN2(g2912), .IN3(n2546), .IN4(g2852), .IN5(
        n2459), .IN6(g2917), .Q(n3328) );
  NOR2X0 U7993 ( .IN1(n3269), .IN2(g904), .QN(g24231) );
  NOR2X0 U7994 ( .IN1(n3261), .IN2(g1249), .QN(g24247) );
  AO21X1 U7995 ( .IN1(g23683), .IN2(n6122), .IN3(n1447), .Q(g24245) );
  AO222X1 U7996 ( .IN1(n2969), .IN2(n3242), .IN3(n2957), .IN4(g1668), .IN5(
        g1636), .IN6(n6098), .Q(g33546) );
  AO222X1 U7997 ( .IN1(n1442), .IN2(g504), .IN3(n1441), .IN4(n2075), .IN5(
        test_so54), .IN6(n5110), .Q(g25610) );
  AO222X1 U7998 ( .IN1(n3091), .IN2(g3352), .IN3(n3092), .IN4(n3093), .IN5(
        g3347), .IN6(n6099), .Q(g33609) );
  NOR2X0 U7999 ( .IN1(g3352), .IN2(n3086), .QN(n3092) );
  AO222X1 U8000 ( .IN1(n3081), .IN2(g3703), .IN3(n3082), .IN4(n3083), .IN5(
        g3698), .IN6(n6099), .Q(g33611) );
  NOR2X0 U8001 ( .IN1(g3703), .IN2(n3075), .QN(n3082) );
  AO222X1 U8002 ( .IN1(n3049), .IN2(g5703), .IN3(n3050), .IN4(n3051), .IN5(
        g5698), .IN6(n6099), .Q(g33620) );
  NOR2X0 U8003 ( .IN1(g5703), .IN2(n3043), .QN(n3050) );
  AO222X1 U8004 ( .IN1(n1305), .IN2(g4975), .IN3(n2758), .IN4(n1607), .IN5(
        g4966), .IN6(n6095), .Q(g34037) );
  INVX0 U8005 ( .IN(n2751), .QN(n1607) );
  NOR2X0 U8006 ( .IN1(g4975), .IN2(n1307), .QN(n2758) );
  AO222X1 U8007 ( .IN1(n3020), .IN2(g6741), .IN3(n3021), .IN4(n3022), .IN5(
        g6736), .IN6(n6100), .Q(g33626) );
  NOR2X0 U8008 ( .IN1(g6741), .IN2(n3014), .QN(n3021) );
  AO222X1 U8009 ( .IN1(n1301), .IN2(g4785), .IN3(n2773), .IN4(n1552), .IN5(
        g4776), .IN6(n6094), .Q(g34029) );
  INVX0 U8010 ( .IN(n2766), .QN(n1552) );
  NOR2X0 U8011 ( .IN1(g4785), .IN2(n1303), .QN(n2773) );
  AO222X1 U8012 ( .IN1(n3057), .IN2(g5357), .IN3(n3058), .IN4(n3059), .IN5(
        g5352), .IN6(n6099), .Q(g33618) );
  NOR2X0 U8013 ( .IN1(g5357), .IN2(n3052), .QN(n3058) );
  AO222X1 U8014 ( .IN1(n3040), .IN2(test_so57), .IN3(n3041), .IN4(n3042), 
        .IN5(test_so50), .IN6(n6099), .Q(g33622) );
  NOR2X0 U8015 ( .IN1(test_so57), .IN2(n3034), .QN(n3041) );
  AO222X1 U8016 ( .IN1(n3072), .IN2(g4054), .IN3(n3073), .IN4(n3074), .IN5(
        g4049), .IN6(n6099), .Q(g33613) );
  NOR2X0 U8017 ( .IN1(g4054), .IN2(n3066), .QN(n3073) );
  AO222X1 U8018 ( .IN1(n3030), .IN2(g6395), .IN3(n3031), .IN4(n3032), .IN5(
        g6390), .IN6(n6100), .Q(g33624) );
  NOR2X0 U8019 ( .IN1(g6395), .IN2(n3024), .QN(n3031) );
  AO222X1 U8020 ( .IN1(n2593), .IN2(n2594), .IN3(n2595), .IN4(g4332), .IN5(
        g4322), .IN6(n6098), .Q(g34455) );
  NOR2X0 U8021 ( .IN1(n5506), .IN2(n2596), .QN(n2593) );
  AO222X1 U8022 ( .IN1(n2899), .IN2(n3183), .IN3(n2887), .IN4(g2070), .IN5(
        g2040), .IN6(n6098), .Q(g33570) );
  AO222X1 U8023 ( .IN1(n2923), .IN2(n3203), .IN3(n2911), .IN4(g1936), .IN5(
        g1906), .IN6(n6098), .Q(g33562) );
  AO222X1 U8024 ( .IN1(n2946), .IN2(n3223), .IN3(n2934), .IN4(g1802), .IN5(
        g1772), .IN6(n6098), .Q(g33554) );
  AO222X1 U8025 ( .IN1(n2853), .IN2(n3143), .IN3(n2840), .IN4(g2361), .IN5(
        g2331), .IN6(n6099), .Q(g33586) );
  AO222X1 U8026 ( .IN1(n2876), .IN2(n3162), .IN3(n2863), .IN4(g2227), .IN5(
        g2197), .IN6(n6098), .Q(g33578) );
  AO222X1 U8027 ( .IN1(g21245), .IN2(n3057), .IN3(n3059), .IN4(n4282), .IN5(
        g5272), .IN6(n6106), .Q(g28093) );
  AO222X1 U8028 ( .IN1(n2753), .IN2(test_so58), .IN3(n1305), .IN4(g4966), 
        .IN5(test_so58), .IN6(n6097), .Q(g34039) );
  NOR2X0 U8029 ( .IN1(n2754), .IN2(n2755), .QN(n2753) );
  AO222X1 U8030 ( .IN1(n2768), .IN2(test_so29), .IN3(n1301), .IN4(g4776), 
        .IN5(test_so29), .IN6(n6095), .Q(g34031) );
  NOR2X0 U8031 ( .IN1(n2769), .IN2(n2770), .QN(n2768) );
  AO222X1 U8032 ( .IN1(n5025), .IN2(g4169), .IN3(n5026), .IN4(n1436), .IN5(
        g4057), .IN6(n6108), .Q(g25687) );
  NOR2X0 U8033 ( .IN1(g4141), .IN2(n4723), .QN(n5025) );
  ISOLANDX1 U8034 ( .D(n4723), .ISO(n5612), .Q(n5026) );
  AO222X1 U8035 ( .IN1(n3940), .IN2(g4169), .IN3(n3941), .IN4(n1436), .IN5(
        g4087), .IN6(n6110), .Q(g30456) );
  ISOLANDX1 U8036 ( .D(n3729), .ISO(n5340), .Q(n3941) );
  NOR2X0 U8037 ( .IN1(g4093), .IN2(n3729), .QN(n3940) );
  AO222X1 U8038 ( .IN1(n1443), .IN2(test_so72), .IN3(n5119), .IN4(g446), .IN5(
        g405), .IN6(n6106), .Q(g25602) );
  AO222X1 U8039 ( .IN1(n1449), .IN2(g392), .IN3(n5252), .IN4(n1448), .IN5(g401), .IN6(n6109), .Q(g24200) );
  NOR2X0 U8040 ( .IN1(g703), .IN2(n5754), .QN(n5252) );
  AO222X1 U8041 ( .IN1(g4035), .IN2(n3072), .IN3(n3074), .IN4(n4343), .IN5(
        g3965), .IN6(n6107), .Q(g28069) );
  AO222X1 U8042 ( .IN1(g3808), .IN2(n3072), .IN3(n4341), .IN4(n3074), .IN5(
        g3813), .IN6(n6107), .Q(g29269) );
  XNOR2X1 U8043 ( .IN1(n4342), .IN2(n4343), .Q(n4341) );
  NAND2X0 U8044 ( .IN1(g3808), .IN2(n4340), .QN(n4342) );
  AO222X1 U8045 ( .IN1(g4826), .IN2(n3030), .IN3(n3032), .IN4(n4237), .IN5(
        g6311), .IN6(n6105), .Q(g28102) );
  AO222X1 U8046 ( .IN1(g6154), .IN2(n3030), .IN3(n4235), .IN4(n3032), .IN5(
        g6159), .IN6(n6108), .Q(g29298) );
  XNOR2X1 U8047 ( .IN1(n4236), .IN2(n4237), .Q(n4235) );
  NAND2X0 U8048 ( .IN1(g6154), .IN2(n4234), .QN(n4236) );
  AO222X1 U8049 ( .IN1(n3732), .IN2(g1367), .IN3(n3733), .IN4(n3658), .IN5(
        g1361), .IN6(n6102), .Q(g31871) );
  ISOLANDX1 U8050 ( .D(n3660), .ISO(g1367), .Q(n3733) );
  NOR2X0 U8051 ( .IN1(n3660), .IN2(n6070), .QN(n3732) );
  AO222X1 U8052 ( .IN1(g4821), .IN2(n3049), .IN3(n3051), .IN4(n4267), .IN5(
        g5619), .IN6(n6106), .Q(g28096) );
  AO222X1 U8053 ( .IN1(n4798), .IN2(n1837), .IN3(n4799), .IN4(n3658), .IN5(
        g1351), .IN6(n6107), .Q(g28059) );
  NOR2X0 U8054 ( .IN1(g1345), .IN2(n1837), .QN(n4799) );
  ISOLANDX1 U8055 ( .D(g1345), .ISO(n6144), .Q(n4798) );
  AO222X1 U8056 ( .IN1(g1636), .IN2(n2957), .IN3(n3250), .IN4(n2972), .IN5(
        test_so75), .IN6(n6098), .Q(g33545) );
  NOR2X0 U8057 ( .IN1(n1289), .IN2(n6067), .QN(n3250) );
  AO222X1 U8058 ( .IN1(n4805), .IN2(n1927), .IN3(n4806), .IN4(n3667), .IN5(
        g1008), .IN6(n6107), .Q(g28057) );
  NOR2X0 U8059 ( .IN1(g1002), .IN2(n1927), .QN(n4806) );
  ISOLANDX1 U8060 ( .D(g1002), .ISO(n6144), .Q(n4805) );
  AO222X1 U8061 ( .IN1(n2599), .IN2(n2598), .IN3(n2600), .IN4(n2591), .IN5(
        g4593), .IN6(n6098), .Q(g34453) );
  NOR2X0 U8062 ( .IN1(n2598), .IN2(n5365), .QN(n2600) );
  NOR2X0 U8063 ( .IN1(g4601), .IN2(n2592), .QN(n2599) );
  AO222X1 U8064 ( .IN1(g5011), .IN2(n3020), .IN3(n3022), .IN4(n4222), .IN5(
        g6657), .IN6(n6110), .Q(g28105) );
  AO222X1 U8065 ( .IN1(n4812), .IN2(n4519), .IN3(n4813), .IN4(n4518), .IN5(
        g822), .IN6(n6107), .Q(g28055) );
  NOR2X0 U8066 ( .IN1(g827), .IN2(n4520), .QN(n4812) );
  NOR2X0 U8067 ( .IN1(n4519), .IN2(n5728), .QN(n4813) );
  AO222X1 U8068 ( .IN1(g3333), .IN2(n3091), .IN3(n3093), .IN4(n4373), .IN5(
        g3263), .IN6(n6107), .Q(g28063) );
  AO222X1 U8069 ( .IN1(n4174), .IN2(g1361), .IN3(n4175), .IN4(n3658), .IN5(
        g1345), .IN6(n6109), .Q(g30343) );
  ISOLANDX1 U8070 ( .D(n3734), .ISO(g1361), .Q(n4175) );
  NOR2X0 U8071 ( .IN1(n3734), .IN2(n6071), .QN(n4174) );
  AO222X1 U8072 ( .IN1(g3684), .IN2(n3081), .IN3(n3083), .IN4(n4358), .IN5(
        g3614), .IN6(n6107), .Q(g28066) );
  AO222X1 U8073 ( .IN1(n4192), .IN2(g1018), .IN3(n4193), .IN4(n3667), .IN5(
        g1002), .IN6(n6108), .Q(g30337) );
  ISOLANDX1 U8074 ( .D(n3739), .ISO(g1018), .Q(n4193) );
  NOR2X0 U8075 ( .IN1(n3739), .IN2(n6071), .QN(n4192) );
  AO222X1 U8076 ( .IN1(n3665), .IN2(g1030), .IN3(n3666), .IN4(n3667), .IN5(
        g1024), .IN6(n6100), .Q(g32983) );
  NOR2X0 U8077 ( .IN1(g1030), .IN2(n1582), .QN(n3666) );
  NOR2X0 U8078 ( .IN1(n3668), .IN2(n6070), .QN(n3665) );
  AO222X1 U8079 ( .IN1(n3656), .IN2(g1373), .IN3(n3657), .IN4(n3658), .IN5(
        g1367), .IN6(n6100), .Q(g32986) );
  NOR2X0 U8080 ( .IN1(g1373), .IN2(n1572), .QN(n3657) );
  NOR2X0 U8081 ( .IN1(n3659), .IN2(n6070), .QN(n3656) );
  AO222X1 U8082 ( .IN1(n2934), .IN2(g1816), .IN3(n2935), .IN4(n2936), .IN5(
        g1802), .IN6(n6101), .Q(g33978) );
  NOR2X0 U8083 ( .IN1(n1356), .IN2(n6065), .QN(n2935) );
  XNOR2X1 U8084 ( .IN1(n2937), .IN2(n2938), .Q(n2936) );
  OA21X1 U8085 ( .IN1(g1728), .IN2(g1802), .IN3(g1816), .Q(n2937) );
  AO222X1 U8086 ( .IN1(g4831), .IN2(n3040), .IN3(n3042), .IN4(n4252), .IN5(
        test_so13), .IN6(n6106), .Q(g28099) );
  AO222X1 U8087 ( .IN1(n3737), .IN2(g1024), .IN3(n3738), .IN4(n3667), .IN5(
        g1018), .IN6(n6102), .Q(g31869) );
  ISOLANDX1 U8088 ( .D(n3669), .ISO(g1024), .Q(n3738) );
  NOR2X0 U8089 ( .IN1(n3669), .IN2(n6070), .QN(n3737) );
  AO222X1 U8090 ( .IN1(g3106), .IN2(n3091), .IN3(n4371), .IN4(n3093), .IN5(
        g3111), .IN6(n6107), .Q(g29257) );
  XNOR2X1 U8091 ( .IN1(n4372), .IN2(n4373), .Q(n4371) );
  NAND2X0 U8092 ( .IN1(g3106), .IN2(n4370), .QN(n4372) );
  AO222X1 U8093 ( .IN1(g5115), .IN2(n3057), .IN3(n4280), .IN4(n3059), .IN5(
        g5120), .IN6(n6107), .Q(g29280) );
  XNOR2X1 U8094 ( .IN1(n4281), .IN2(n4282), .Q(n4280) );
  NAND2X0 U8095 ( .IN1(g5115), .IN2(n4279), .QN(n4281) );
  AO222X1 U8096 ( .IN1(n4863), .IN2(n4861), .IN3(n4866), .IN4(g4438), .IN5(
        test_so47), .IN6(n6109), .Q(g26954) );
  AO222X1 U8097 ( .IN1(g2779), .IN2(n4888), .IN3(n4889), .IN4(n5834), .IN5(
        g2767), .IN6(n6110), .Q(g26928) );
  AO222X1 U8098 ( .IN1(n4721), .IN2(n4716), .IN3(n4717), .IN4(g4119), .IN5(
        g4116), .IN6(n6106), .Q(g28073) );
  NOR2X0 U8099 ( .IN1(n4716), .IN2(n6068), .QN(n4717) );
  AND3X1 U8100 ( .IN1(g4057), .IN2(n5416), .IN3(n4722), .Q(n4716) );
  AO222X1 U8101 ( .IN1(n4888), .IN2(g2827), .IN3(n4889), .IN4(n5835), .IN5(
        test_so37), .IN6(n6109), .Q(g26934) );
  AO222X1 U8102 ( .IN1(n2558), .IN2(g4854), .IN3(n2559), .IN4(g4859), .IN5(
        g4854), .IN6(n6097), .Q(g34468) );
  NOR2X0 U8103 ( .IN1(n2560), .IN2(n2561), .QN(n2558) );
  AO222X1 U8104 ( .IN1(n2605), .IN2(n2594), .IN3(n2606), .IN4(n2595), .IN5(
        g4311), .IN6(n6098), .Q(g34450) );
  NOR2X0 U8105 ( .IN1(n2594), .IN2(n5506), .QN(n2606) );
  NOR2X0 U8106 ( .IN1(g4322), .IN2(n2596), .QN(n2605) );
  AO222X1 U8107 ( .IN1(g5462), .IN2(n3049), .IN3(n4265), .IN4(n3051), .IN5(
        g5467), .IN6(n6107), .Q(g29286) );
  XNOR2X1 U8108 ( .IN1(n4266), .IN2(n4267), .Q(n4265) );
  NAND2X0 U8109 ( .IN1(g5462), .IN2(n4264), .QN(n4266) );
  AO222X1 U8110 ( .IN1(n4522), .IN2(n4523), .IN3(n4524), .IN4(test_so70), 
        .IN5(g676), .IN6(n6106), .Q(g29227) );
  NOR2X0 U8111 ( .IN1(test_so70), .IN2(n4527), .QN(n4522) );
  ISOLANDX1 U8112 ( .D(n4525), .ISO(n4523), .Q(n4524) );
  ISOLANDX1 U8113 ( .D(n4526), .ISO(n5751), .Q(n4523) );
  AO222X1 U8114 ( .IN1(g2767), .IN2(n4888), .IN3(n4889), .IN4(n5836), .IN5(
        g2763), .IN6(n6110), .Q(g26927) );
  AO222X1 U8115 ( .IN1(g2791), .IN2(n4888), .IN3(n4889), .IN4(n5837), .IN5(
        g2779), .IN6(n6109), .Q(g26929) );
  AO222X1 U8116 ( .IN1(n4888), .IN2(g2795), .IN3(n4889), .IN4(n5838), .IN5(
        g2791), .IN6(n6109), .Q(g26930) );
  AO222X1 U8117 ( .IN1(g2799), .IN2(n4888), .IN3(n4889), .IN4(n5839), .IN5(
        g20654), .IN6(n6109), .Q(g26931) );
  AO222X1 U8118 ( .IN1(g6500), .IN2(n3020), .IN3(n4220), .IN4(n3022), .IN5(
        g6505), .IN6(n6108), .Q(g29304) );
  XNOR2X1 U8119 ( .IN1(n4221), .IN2(n4222), .Q(n4220) );
  NAND2X0 U8120 ( .IN1(g6500), .IN2(n4219), .QN(n4221) );
  AO222X1 U8121 ( .IN1(n4721), .IN2(n4718), .IN3(n4719), .IN4(g4116), .IN5(
        g4112), .IN6(n6106), .Q(g28072) );
  NOR2X0 U8122 ( .IN1(n4718), .IN2(n6068), .QN(n4719) );
  AND3X1 U8123 ( .IN1(g4064), .IN2(n5711), .IN3(n4722), .Q(n4718) );
  AO222X1 U8124 ( .IN1(n2568), .IN2(g4664), .IN3(n2569), .IN4(g4669), .IN5(
        g4664), .IN6(n6098), .Q(g34464) );
  NOR2X0 U8125 ( .IN1(n2570), .IN2(n2571), .QN(n2568) );
  AO222X1 U8126 ( .IN1(test_so37), .IN2(n4888), .IN3(n4889), .IN4(n5840), 
        .IN5(g2811), .IN6(n6109), .Q(g26933) );
  AO222X1 U8127 ( .IN1(g2811), .IN2(n4888), .IN3(n4889), .IN4(n5841), .IN5(
        g2799), .IN6(n6109), .Q(g26932) );
  AO222X1 U8128 ( .IN1(g5808), .IN2(n3040), .IN3(n4250), .IN4(n3042), .IN5(
        g5813), .IN6(n6108), .Q(g29292) );
  XNOR2X1 U8129 ( .IN1(n4251), .IN2(n4252), .Q(n4250) );
  NAND2X0 U8130 ( .IN1(g5808), .IN2(n4249), .QN(n4251) );
  AO222X1 U8131 ( .IN1(n3699), .IN2(n3700), .IN3(n3701), .IN4(n1399), .IN5(
        g5016), .IN6(n6101), .Q(g31902) );
  NOR2X0 U8132 ( .IN1(n3700), .IN2(n5601), .QN(n3701) );
  OA22X1 U8133 ( .IN1(n5369), .IN2(g5062), .IN3(g5016), .IN4(g5022), .Q(n3700)
         );
  NOR2X0 U8134 ( .IN1(g5029), .IN2(n6070), .QN(n3699) );
  AO222X1 U8135 ( .IN1(n3713), .IN2(n6167), .IN3(n3714), .IN4(n3715), .IN5(
        g5033), .IN6(n6101), .Q(g31899) );
  NOR2X0 U8136 ( .IN1(g5037), .IN2(n3715), .QN(n3713) );
  NOR2X0 U8137 ( .IN1(n5611), .IN2(n3451), .QN(n3714) );
  AOI21X1 U8138 ( .IN1(g5033), .IN2(n1874), .IN3(n3688), .QN(n3715) );
  AO222X1 U8139 ( .IN1(test_so4), .IN2(n3081), .IN3(n4356), .IN4(n3083), .IN5(
        g3462), .IN6(n6107), .Q(g29263) );
  XNOR2X1 U8140 ( .IN1(n4357), .IN2(n4358), .Q(n4356) );
  NAND2X0 U8141 ( .IN1(test_so4), .IN2(n4355), .QN(n4357) );
  AO222X1 U8142 ( .IN1(n3448), .IN2(n6166), .IN3(n3449), .IN4(n3450), .IN5(
        g5052), .IN6(n6089), .Q(g33046) );
  NOR2X0 U8143 ( .IN1(g5057), .IN2(n3450), .QN(n3448) );
  NOR2X0 U8144 ( .IN1(n5615), .IN2(n3451), .QN(n3449) );
  AOI21X1 U8145 ( .IN1(g5052), .IN2(n1822), .IN3(n3452), .QN(n3450) );
  AO222X1 U8146 ( .IN1(n2576), .IN2(n2573), .IN3(n2577), .IN4(n2569), .IN5(
        test_so19), .IN6(n6098), .Q(g34461) );
  ISOLANDX1 U8147 ( .D(g4659), .ISO(n2573), .Q(n2577) );
  NOR2X0 U8148 ( .IN1(g4659), .IN2(n2570), .QN(n2576) );
  AO222X1 U8149 ( .IN1(n3716), .IN2(n3717), .IN3(n3718), .IN4(n1399), .IN5(
        g5022), .IN6(n6101), .Q(g31898) );
  NOR2X0 U8150 ( .IN1(g5016), .IN2(n3717), .QN(n3718) );
  NOR2X0 U8151 ( .IN1(g5062), .IN2(g5022), .QN(n3717) );
  NOR2X0 U8152 ( .IN1(n6083), .IN2(n5369), .QN(n3716) );
  AO222X1 U8153 ( .IN1(n2425), .IN2(n5292), .IN3(n2484), .IN4(n2404), .IN5(
        g785), .IN6(n6095), .Q(g34791) );
  NOR2X0 U8154 ( .IN1(n2425), .IN2(n5292), .QN(n2484) );
  AO222X1 U8155 ( .IN1(g872), .IN2(n4944), .IN3(n4945), .IN4(g446), .IN5(g246), 
        .IN6(n6114), .Q(g26908) );
  AO222X1 U8156 ( .IN1(g650), .IN2(n1421), .IN3(n4816), .IN4(g681), .IN5(
        test_so87), .IN6(n6108), .Q(g28049) );
  AO222X1 U8157 ( .IN1(n2485), .IN2(n5293), .IN3(n2506), .IN4(n2404), .IN5(
        g781), .IN6(n6094), .Q(g34725) );
  NOR2X0 U8158 ( .IN1(n2485), .IN2(n5293), .QN(n2506) );
  AO222X1 U8159 ( .IN1(n2507), .IN2(n5551), .IN3(n2553), .IN4(n2404), .IN5(
        g776), .IN6(n6097), .Q(g34600) );
  NOR2X0 U8160 ( .IN1(n2507), .IN2(n5551), .QN(n2553) );
  AO222X1 U8161 ( .IN1(n2554), .IN2(n5330), .IN3(n2646), .IN4(n2404), .IN5(
        g772), .IN6(n6091), .Q(g34439) );
  NOR2X0 U8162 ( .IN1(n2554), .IN2(n5330), .QN(n2646) );
  AO222X1 U8163 ( .IN1(g475), .IN2(n1449), .IN3(n1448), .IN4(g246), .IN5(g424), 
        .IN6(n6109), .Q(g24208) );
  AO222X1 U8164 ( .IN1(n2566), .IN2(n2563), .IN3(n2567), .IN4(n2559), .IN5(
        g4843), .IN6(n6097), .Q(g34465) );
  ISOLANDX1 U8165 ( .D(g4849), .ISO(n2563), .Q(n2567) );
  NOR2X0 U8166 ( .IN1(g4849), .IN2(n2560), .QN(n2566) );
  AO222X1 U8167 ( .IN1(n3272), .IN2(n5331), .IN3(n3681), .IN4(n2404), .IN5(
        test_so2), .IN6(n6100), .Q(g32979) );
  NOR2X0 U8168 ( .IN1(n3272), .IN2(n5331), .QN(n3681) );
  AO222X1 U8169 ( .IN1(test_so23), .IN2(n1449), .IN3(n1448), .IN4(g269), .IN5(
        g437), .IN6(n6109), .Q(g24205) );
  AO222X1 U8170 ( .IN1(n3743), .IN2(n5470), .IN3(n4197), .IN4(n2404), .IN5(
        test_so60), .IN6(n6108), .Q(g30335) );
  NOR2X0 U8171 ( .IN1(n3743), .IN2(n5470), .QN(n4197) );
  AO222X1 U8172 ( .IN1(n2980), .IN2(n5332), .IN3(n3271), .IN4(n2404), .IN5(
        g758), .IN6(n6097), .Q(g33539) );
  NOR2X0 U8173 ( .IN1(n2980), .IN2(n5332), .QN(n3271) );
  AO222X1 U8174 ( .IN1(n2704), .IN2(n5333), .IN3(n2979), .IN4(n2404), .IN5(
        g763), .IN6(n6100), .Q(g33965) );
  NOR2X0 U8175 ( .IN1(n2704), .IN2(n5333), .QN(n2979) );
  AO222X1 U8176 ( .IN1(n2647), .IN2(n5334), .IN3(n2703), .IN4(n2404), .IN5(
        g767), .IN6(n6093), .Q(g34252) );
  NOR2X0 U8177 ( .IN1(n2647), .IN2(n5334), .QN(n2703) );
  AO222X1 U8178 ( .IN1(n3682), .IN2(n5471), .IN3(n3742), .IN4(n2404), .IN5(
        g744), .IN6(n6102), .Q(g31867) );
  NOR2X0 U8179 ( .IN1(n3682), .IN2(n5471), .QN(n3742) );
  AO222X1 U8180 ( .IN1(n5019), .IN2(g5077), .IN3(n5020), .IN4(n1435), .IN5(
        g5080), .IN6(n5021), .Q(g25696) );
  OA21X1 U8181 ( .IN1(g5069), .IN2(n5455), .IN3(n5893), .Q(n5020) );
  INVX0 U8182 ( .IN(n5021), .QN(n1435) );
  NAND2X0 U8183 ( .IN1(n6210), .IN2(n5681), .QN(n5021) );
  AO222X1 U8184 ( .IN1(n4937), .IN2(g1046), .IN3(n4938), .IN4(n4939), .IN5(
        g1041), .IN6(n6110), .Q(g26913) );
  ISOLANDX1 U8185 ( .D(n4940), .ISO(g1046), .Q(n4938) );
  NOR2X0 U8186 ( .IN1(n4940), .IN2(n6066), .QN(n4937) );
  OA21X1 U8187 ( .IN1(n5321), .IN2(g1041), .IN3(n1928), .Q(n4940) );
  AO222X1 U8188 ( .IN1(n5085), .IN2(g1041), .IN3(n5086), .IN4(n4939), .IN5(
        g1036), .IN6(n6106), .Q(g25624) );
  NOR2X0 U8189 ( .IN1(g1041), .IN2(n5087), .QN(n5086) );
  NOR2X0 U8190 ( .IN1(n1928), .IN2(n6078), .QN(n5085) );
  AO222X1 U8191 ( .IN1(n4912), .IN2(g1389), .IN3(n4913), .IN4(n4914), .IN5(
        g1384), .IN6(n6115), .Q(g26920) );
  ISOLANDX1 U8192 ( .D(n4915), .ISO(g1389), .Q(n4913) );
  NOR2X0 U8193 ( .IN1(n4915), .IN2(n6066), .QN(n4912) );
  OA21X1 U8194 ( .IN1(n5322), .IN2(g1384), .IN3(n1574), .Q(n4915) );
  AO222X1 U8195 ( .IN1(n4528), .IN2(n4526), .IN3(n4529), .IN4(n4525), .IN5(
        g671), .IN6(n6105), .Q(g29226) );
  NOR2X0 U8196 ( .IN1(n4526), .IN2(n5751), .QN(n4529) );
  NOR2X0 U8197 ( .IN1(g676), .IN2(n4527), .QN(n4528) );
  AO222X1 U8198 ( .IN1(n5061), .IN2(g1384), .IN3(n5062), .IN4(n4914), .IN5(
        g1379), .IN6(n6107), .Q(g25633) );
  NOR2X0 U8199 ( .IN1(g1384), .IN2(n5063), .QN(n5062) );
  NOR2X0 U8200 ( .IN1(n1574), .IN2(n6079), .QN(n5061) );
  AO222X1 U8201 ( .IN1(g14201), .IN2(n4944), .IN3(n4945), .IN4(g255), .IN5(
        g225), .IN6(n6110), .Q(g26902) );
  AO222X1 U8202 ( .IN1(g14096), .IN2(n4944), .IN3(n4945), .IN4(g262), .IN5(
        g232), .IN6(n6110), .Q(g26904) );
  AO222X1 U8203 ( .IN1(g14217), .IN2(n4944), .IN3(n4945), .IN4(g232), .IN5(
        g255), .IN6(n6110), .Q(g26903) );
  AO222X1 U8204 ( .IN1(g14125), .IN2(n4944), .IN3(n4945), .IN4(g239), .IN5(
        g262), .IN6(n6110), .Q(g26905) );
  AO222X1 U8205 ( .IN1(g14147), .IN2(n4944), .IN3(n4945), .IN4(g269), .IN5(
        g239), .IN6(n6110), .Q(g26906) );
  AO222X1 U8206 ( .IN1(g14189), .IN2(n4944), .IN3(n4945), .IN4(g225), .IN5(
        g872), .IN6(n6110), .Q(g26901) );
  AO222X1 U8207 ( .IN1(g14167), .IN2(n4944), .IN3(n4945), .IN4(g246), .IN5(
        g269), .IN6(n6114), .Q(g26907) );
  AO222X1 U8208 ( .IN1(n4721), .IN2(n4714), .IN3(n4715), .IN4(g4122), .IN5(
        g4119), .IN6(n6106), .Q(g28074) );
  NOR2X0 U8209 ( .IN1(n4714), .IN2(n6068), .QN(n4715) );
  ISOLANDX1 U8210 ( .D(n4722), .ISO(n4723), .Q(n4714) );
  AO222X1 U8211 ( .IN1(n1871), .IN2(n5730), .IN3(n3260), .IN4(g1274), .IN5(
        g1270), .IN6(n6097), .Q(g33542) );
  NOR2X0 U8212 ( .IN1(n1871), .IN2(n3261), .QN(n3260) );
  INVX0 U8213 ( .IN(n3262), .QN(n1871) );
  AO222X1 U8214 ( .IN1(n1604), .IN2(n5731), .IN3(n3268), .IN4(g930), .IN5(g925), .IN6(n6097), .Q(g33540) );
  NOR2X0 U8215 ( .IN1(n1604), .IN2(n3269), .QN(n3268) );
  INVX0 U8216 ( .IN(n3270), .QN(n1604) );
  AO222X1 U8217 ( .IN1(n5078), .IN2(n1694), .IN3(n5079), .IN4(g962), .IN5(
        g1178), .IN6(n6106), .Q(g25627) );
  OA21X1 U8218 ( .IN1(n3215), .IN2(n5304), .IN3(n6367), .Q(n5079) );
  AO222X1 U8219 ( .IN1(n2589), .IN2(n2590), .IN3(n2591), .IN4(g4616), .IN5(
        g4608), .IN6(n6098), .Q(g34456) );
  NOR2X0 U8220 ( .IN1(n5274), .IN2(n2592), .QN(n2589) );
  AO222X1 U8221 ( .IN1(n4515), .IN2(n4516), .IN3(n4517), .IN4(g723), .IN5(g827), .IN6(n6106), .Q(g29229) );
  NOR2X0 U8222 ( .IN1(g723), .IN2(n4520), .QN(n4515) );
  ISOLANDX1 U8223 ( .D(n4518), .ISO(n4516), .Q(n4517) );
  ISOLANDX1 U8224 ( .D(n4519), .ISO(n5728), .Q(n4516) );
  AO222X1 U8225 ( .IN1(n2710), .IN2(n5843), .IN3(n2711), .IN4(g160), .IN5(g157), .IN6(n6097), .Q(g34249) );
  NOR2X0 U8226 ( .IN1(n2710), .IN2(n2712), .QN(n2711) );
  AO222X1 U8227 ( .IN1(n2707), .IN2(n5724), .IN3(n2708), .IN4(g142), .IN5(g298), .IN6(n6095), .Q(g34250) );
  NOR2X0 U8228 ( .IN1(n2707), .IN2(n2709), .QN(n2708) );
  AO222X1 U8229 ( .IN1(n4177), .IN2(n1445), .IN3(n3736), .IN4(n5553), .IN5(
        g1256), .IN6(n6109), .Q(g30342) );
  NOR2X0 U8230 ( .IN1(n3736), .IN2(n5553), .QN(n4177) );
  AO222X1 U8231 ( .IN1(n3663), .IN2(n1445), .IN3(n3662), .IN4(n5716), .IN5(
        g1263), .IN6(n6100), .Q(g32984) );
  NOR2X0 U8232 ( .IN1(n3662), .IN2(n5716), .QN(n3663) );
  AO222X1 U8233 ( .IN1(n4803), .IN2(n1445), .IN3(n4490), .IN4(n5554), .IN5(
        test_so77), .IN6(n6107), .Q(g28058) );
  NOR2X0 U8234 ( .IN1(n4490), .IN2(n5554), .QN(n4803) );
  AO222X1 U8235 ( .IN1(n4973), .IN2(n1540), .IN3(n4974), .IN4(g336), .IN5(g311), .IN6(n6109), .Q(g26886) );
  NOR2X0 U8236 ( .IN1(n6083), .IN2(n1540), .QN(n4974) );
  AO222X1 U8237 ( .IN1(g460), .IN2(n1443), .IN3(n5119), .IN4(g246), .IN5(g168), 
        .IN6(n6106), .Q(g25605) );
  AO222X1 U8238 ( .IN1(n1279), .IN2(n3493), .IN3(n3494), .IN4(g25648), .IN5(
        g3171), .IN6(n6101), .Q(g33024) );
  NAND2X0 U8239 ( .IN1(n3495), .IN2(n3496), .QN(n3493) );
  AO222X1 U8240 ( .IN1(n3671), .IN2(n5725), .IN3(n3672), .IN4(n1447), .IN5(
        g918), .IN6(n6100), .Q(g32981) );
  NOR2X0 U8241 ( .IN1(n3671), .IN2(n5725), .QN(n3672) );
  AO222X1 U8242 ( .IN1(n2756), .IN2(n1306), .IN3(n2757), .IN4(test_so58), 
        .IN5(g4983), .IN6(n6097), .Q(g34038) );
  NOR2X0 U8243 ( .IN1(test_so58), .IN2(n2754), .QN(n2756) );
  NOR2X0 U8244 ( .IN1(n1608), .IN2(n2748), .QN(n2757) );
  AO222X1 U8245 ( .IN1(n2771), .IN2(n1302), .IN3(n2772), .IN4(test_so29), 
        .IN5(g4793), .IN6(n6094), .Q(g34030) );
  NOR2X0 U8246 ( .IN1(test_so29), .IN2(n2769), .QN(n2771) );
  NOR2X0 U8247 ( .IN1(n1727), .IN2(n2763), .QN(n2772) );
  AO222X1 U8248 ( .IN1(n4514), .IN2(n5555), .IN3(n4810), .IN4(n1447), .IN5(
        g936), .IN6(n6107), .Q(g28056) );
  NOR2X0 U8249 ( .IN1(n4514), .IN2(n5555), .QN(n4810) );
  AO222X1 U8250 ( .IN1(n4804), .IN2(n5556), .IN3(n4916), .IN4(n1445), .IN5(
        g1266), .IN6(n6115), .Q(g26919) );
  NOR2X0 U8251 ( .IN1(n4804), .IN2(n5556), .QN(n4916) );
  AO222X1 U8252 ( .IN1(n4811), .IN2(n5557), .IN3(n4941), .IN4(n1447), .IN5(
        g921), .IN6(n6115), .Q(g26912) );
  NOR2X0 U8253 ( .IN1(n4811), .IN2(n5557), .QN(n4941) );
  AO222X1 U8254 ( .IN1(n2830), .IN2(n1295), .IN3(n2817), .IN4(g2495), .IN5(
        g2465), .IN6(n6099), .Q(g33594) );
  AO222X1 U8255 ( .IN1(n3673), .IN2(n5673), .IN3(n3740), .IN4(n1447), .IN5(
        g914), .IN6(n6102), .Q(g31868) );
  NOR2X0 U8256 ( .IN1(n3673), .IN2(n5673), .QN(n3740) );
  AO222X1 U8257 ( .IN1(n2806), .IN2(n1296), .IN3(n2793), .IN4(g2629), .IN5(
        g2599), .IN6(n6099), .Q(g33602) );
  AO222X1 U8258 ( .IN1(n3664), .IN2(n5674), .IN3(n3735), .IN4(n1445), .IN5(
        g1259), .IN6(n6102), .Q(g31870) );
  NOR2X0 U8259 ( .IN1(n3664), .IN2(n5674), .QN(n3735) );
  AO222X1 U8260 ( .IN1(n4178), .IN2(n5558), .IN3(n4489), .IN4(n1445), .IN5(
        g1252), .IN6(n6106), .Q(g29235) );
  NOR2X0 U8261 ( .IN1(n4178), .IN2(n5558), .QN(n4489) );
  AO222X1 U8262 ( .IN1(n4196), .IN2(n5559), .IN3(n4513), .IN4(n1447), .IN5(
        g907), .IN6(n6106), .Q(g29230) );
  NOR2X0 U8263 ( .IN1(n4196), .IN2(n5559), .QN(n4513) );
  AO222X1 U8264 ( .IN1(n3741), .IN2(n5560), .IN3(n4195), .IN4(n1447), .IN5(
        g911), .IN6(n6108), .Q(g30336) );
  NOR2X0 U8265 ( .IN1(n3741), .IN2(n5560), .QN(n4195) );
  AO222X1 U8266 ( .IN1(n3687), .IN2(n5561), .IN3(n3749), .IN4(n1411), .IN5(
        test_so73), .IN6(n6102), .Q(g31864) );
  NOR2X0 U8267 ( .IN1(n3687), .IN2(n5561), .QN(n3749) );
  AO222X1 U8268 ( .IN1(n2989), .IN2(n5675), .IN3(n2990), .IN4(n1422), .IN5(
        g294), .IN6(n6100), .Q(g33961) );
  NOR2X0 U8269 ( .IN1(n2989), .IN2(n5675), .QN(n2990) );
  AO222X1 U8270 ( .IN1(n3281), .IN2(n5676), .IN3(n3686), .IN4(n1411), .IN5(
        g164), .IN6(n6101), .Q(g32976) );
  NOR2X0 U8271 ( .IN1(n3281), .IN2(n5676), .QN(n3686) );
  AO222X1 U8272 ( .IN1(n3277), .IN2(n5677), .IN3(n3280), .IN4(n1411), .IN5(
        g150), .IN6(n6097), .Q(g33534) );
  NOR2X0 U8273 ( .IN1(n3277), .IN2(n5677), .QN(n3280) );
  AO222X1 U8274 ( .IN1(n2991), .IN2(n5678), .IN3(n2992), .IN4(n1411), .IN5(
        g153), .IN6(n6100), .Q(g33960) );
  NOR2X0 U8275 ( .IN1(n2991), .IN2(n5678), .QN(n2992) );
  AO222X1 U8276 ( .IN1(n3279), .IN2(n5679), .IN3(n3685), .IN4(n1422), .IN5(
        test_so51), .IN6(n6101), .Q(g32977) );
  NOR2X0 U8277 ( .IN1(n3279), .IN2(n5679), .QN(n3685) );
  AO222X1 U8278 ( .IN1(n3276), .IN2(n5680), .IN3(n3278), .IN4(n1422), .IN5(
        g291), .IN6(n6097), .Q(g33535) );
  NOR2X0 U8279 ( .IN1(n3276), .IN2(n5680), .QN(n3278) );
  AO222X1 U8280 ( .IN1(g686), .IN2(n1442), .IN3(n5111), .IN4(n2075), .IN5(g691), .IN6(n6105), .Q(g25614) );
  ISOLANDX1 U8281 ( .D(n4819), .ISO(n6144), .Q(n5111) );
  AO222X1 U8282 ( .IN1(g1740), .IN2(n1357), .IN3(n2932), .IN4(n1358), .IN5(
        g1821), .IN6(n6101), .Q(g33979) );
  NOR2X0 U8283 ( .IN1(n2933), .IN2(n6065), .QN(n2932) );
  AO222X1 U8284 ( .IN1(g1874), .IN2(n1366), .IN3(n2909), .IN4(n1367), .IN5(
        g1955), .IN6(n6102), .Q(g33986) );
  NOR2X0 U8285 ( .IN1(n2910), .IN2(n6065), .QN(n2909) );
  AO222X1 U8286 ( .IN1(g2165), .IN2(n1310), .IN3(n2861), .IN4(n1311), .IN5(
        g2246), .IN6(n6091), .Q(g34000) );
  NOR2X0 U8287 ( .IN1(n2862), .IN2(n6064), .QN(n2861) );
  AO222X1 U8288 ( .IN1(g2567), .IN2(n1334), .IN3(n2791), .IN4(n1335), .IN5(
        g2648), .IN6(n6093), .Q(g34021) );
  NOR2X0 U8289 ( .IN1(n2792), .IN2(n6063), .QN(n2791) );
  AO222X1 U8290 ( .IN1(g2433), .IN2(n1326), .IN3(n2815), .IN4(n1327), .IN5(
        g2514), .IN6(n6093), .Q(g34014) );
  NOR2X0 U8291 ( .IN1(n2816), .IN2(n6064), .QN(n2815) );
  AO222X1 U8292 ( .IN1(g2008), .IN2(n1375), .IN3(n2885), .IN4(n1376), .IN5(
        g2089), .IN6(n6104), .Q(g33993) );
  NOR2X0 U8293 ( .IN1(n2886), .IN2(n6065), .QN(n2885) );
  AO222X1 U8294 ( .IN1(g1604), .IN2(n1348), .IN3(n2955), .IN4(n1349), .IN5(
        g1687), .IN6(n6101), .Q(g33972) );
  NOR2X0 U8295 ( .IN1(n2956), .IN2(n6065), .QN(n2955) );
  AO222X1 U8296 ( .IN1(g2299), .IN2(n1318), .IN3(n2838), .IN4(n1319), .IN5(
        g2380), .IN6(n6092), .Q(g34007) );
  NOR2X0 U8297 ( .IN1(n2839), .IN2(n6064), .QN(n2838) );
  NOR2X0 U8298 ( .IN1(g6203), .IN2(n3411), .QN(g30522) );
  NOR2X0 U8299 ( .IN1(g3857), .IN2(n3476), .QN(g30435) );
  NOR2X0 U8300 ( .IN1(g5857), .IN2(n3421), .QN(g30501) );
  NOR2X0 U8301 ( .IN1(g6549), .IN2(n3401), .QN(g30543) );
  NOR2X0 U8302 ( .IN1(g5164), .IN2(n3441), .QN(g30459) );
  NOR2X0 U8303 ( .IN1(g5511), .IN2(n3431), .QN(g30480) );
  NOR2X0 U8304 ( .IN1(g3506), .IN2(n3486), .QN(g30414) );
  AO22X1 U8305 ( .IN1(g316), .IN2(n6269), .IN3(g21176), .IN4(n6137), .Q(g26888) );
  AO22X1 U8306 ( .IN1(test_so76), .IN2(n6125), .IN3(g20901), .IN4(n6282), .Q(
        g24242) );
  ISOLANDX1 U8307 ( .D(g21176), .ISO(n6145), .Q(g26900) );
  AND2X1 U8308 ( .IN1(n5979), .IN2(n5980), .Q(n2983) );
  AO221X1 U8309 ( .IN1(n5962), .IN2(g269), .IN3(n6018), .IN4(g262), .IN5(n6016), .Q(n5979) );
  AO21X1 U8310 ( .IN1(n5962), .IN2(g255), .IN3(n1492), .Q(n5980) );
  NOR4X0 U8311 ( .IN1(n5152), .IN2(g17607), .IN3(g13068), .IN4(g17646), .QN(
        g24344) );
  AO221X1 U8312 ( .IN1(g17739), .IN2(n5698), .IN3(g14738), .IN4(n5432), .IN5(
        n6083), .Q(n5152) );
  OA21X1 U8313 ( .IN1(g817), .IN2(n6118), .IN3(n4545), .Q(n5099) );
  AO21X1 U8314 ( .IN1(g20049), .IN2(n6121), .IN3(g29277), .Q(g29276) );
  NAND2X0 U8315 ( .IN1(g3466), .IN2(n6150), .QN(n2475) );
  NAND2X0 U8316 ( .IN1(n3177), .IN2(DFF_1092_n1), .QN(n4473) );
  NAND2X0 U8317 ( .IN1(n3254), .IN2(DFF_24_n1), .QN(n4497) );
  NAND2X0 U8318 ( .IN1(g3817), .IN2(n6152), .QN(n2478) );
  AO22X1 U8319 ( .IN1(g2719), .IN2(n6130), .IN3(n3730), .IN4(n4891), .Q(g26926) );
  XNOR2X1 U8320 ( .IN1(g2724), .IN2(n4052), .Q(n4891) );
  NOR2X0 U8321 ( .IN1(n6081), .IN2(g4258), .QN(g21893) );
  AO222X1 U8322 ( .IN1(n2616), .IN2(g2775), .IN3(n2633), .IN4(n2618), .IN5(
        g2783), .IN6(n6102), .Q(g34443) );
  NOR2X0 U8323 ( .IN1(n2629), .IN2(n2634), .QN(n2633) );
  OA21X1 U8324 ( .IN1(g2779), .IN2(n6118), .IN3(n2615), .Q(n2634) );
  AO222X1 U8325 ( .IN1(n2624), .IN2(g2803), .IN3(n2625), .IN4(n2626), .IN5(
        g2807), .IN6(n6101), .Q(g34445) );
  NOR2X0 U8326 ( .IN1(n2613), .IN2(n2627), .QN(n2625) );
  OA21X1 U8327 ( .IN1(g2799), .IN2(n6118), .IN3(n2615), .Q(n2627) );
  AO222X1 U8328 ( .IN1(n2610), .IN2(g2787), .IN3(n2628), .IN4(n2612), .IN5(
        g2795), .IN6(n6101), .Q(g34444) );
  NOR2X0 U8329 ( .IN1(n2629), .IN2(n2630), .QN(n2628) );
  OA21X1 U8330 ( .IN1(g2795), .IN2(n6118), .IN3(n2615), .Q(n2630) );
  AO222X1 U8331 ( .IN1(n2620), .IN2(g2783), .IN3(n2635), .IN4(n2622), .IN5(
        g2787), .IN6(n6104), .Q(g34442) );
  NOR2X0 U8332 ( .IN1(n2629), .IN2(n2636), .QN(n2635) );
  OA21X1 U8333 ( .IN1(g2791), .IN2(n6118), .IN3(n2615), .Q(n2636) );
  AO222X1 U8334 ( .IN1(n2620), .IN2(g2815), .IN3(n2621), .IN4(n2622), .IN5(
        g2819), .IN6(n6101), .Q(g34446) );
  NOR2X0 U8335 ( .IN1(n2613), .IN2(n2623), .QN(n2621) );
  OA21X1 U8336 ( .IN1(test_so37), .IN2(n6118), .IN3(n2615), .Q(n2623) );
  AO222X1 U8337 ( .IN1(n2616), .IN2(g2807), .IN3(n2617), .IN4(n2618), .IN5(
        g2815), .IN6(n6099), .Q(g34447) );
  NOR2X0 U8338 ( .IN1(n2613), .IN2(n2619), .QN(n2617) );
  OA21X1 U8339 ( .IN1(g2811), .IN2(n6118), .IN3(n2615), .Q(n2619) );
  AO222X1 U8340 ( .IN1(n2610), .IN2(g2819), .IN3(n2611), .IN4(n2612), .IN5(
        g2827), .IN6(n6099), .Q(g34448) );
  NOR2X0 U8341 ( .IN1(n2613), .IN2(n2614), .QN(n2611) );
  OA21X1 U8342 ( .IN1(g2827), .IN2(n6118), .IN3(n2615), .Q(n2614) );
  AO222X1 U8343 ( .IN1(n2624), .IN2(g2771), .IN3(n2638), .IN4(n2626), .IN5(
        g2775), .IN6(n6090), .Q(g34441) );
  NOR2X0 U8344 ( .IN1(n2629), .IN2(n2639), .QN(n2638) );
  OA21X1 U8345 ( .IN1(g2767), .IN2(n6118), .IN3(n2615), .Q(n2639) );
  AO22X1 U8346 ( .IN1(g854), .IN2(n4545), .IN3(n1449), .IN4(g847), .Q(g24216)
         );
  AO22X1 U8347 ( .IN1(g837), .IN2(n5240), .IN3(g703), .IN4(n5241), .Q(g24215)
         );
  NAND2X0 U8348 ( .IN1(n4545), .IN2(n5242), .QN(n5240) );
  AO21X1 U8349 ( .IN1(n4953), .IN2(n5562), .IN3(n6138), .Q(n5241) );
  NAND3X0 U8350 ( .IN1(n5243), .IN2(n5244), .IN3(n6324), .QN(n5242) );
  AO22X1 U8351 ( .IN1(g411), .IN2(n4545), .IN3(n1449), .IN4(g424), .Q(g24202)
         );
  AO22X1 U8352 ( .IN1(test_so23), .IN2(n4545), .IN3(g429), .IN4(n1449), .Q(
        g24204) );
  AO22X1 U8353 ( .IN1(g392), .IN2(n4545), .IN3(n1449), .IN4(g405), .Q(g24201)
         );
  AO22X1 U8354 ( .IN1(g475), .IN2(n4545), .IN3(g441), .IN4(n1449), .Q(g24207)
         );
  AO22X1 U8355 ( .IN1(g429), .IN2(n4545), .IN3(n1449), .IN4(g401), .Q(g24203)
         );
  AO22X1 U8356 ( .IN1(g441), .IN2(n4545), .IN3(n1449), .IN4(g437), .Q(g24206)
         );
  AO22X1 U8357 ( .IN1(g21893), .IN2(g4264), .IN3(g4258), .IN4(n5263), .Q(
        g21894) );
  NAND2X0 U8358 ( .IN1(g4264), .IN2(n6175), .QN(n5263) );
  AO22X1 U8359 ( .IN1(n3091), .IN2(g4939), .IN3(n4683), .IN4(n1701), .Q(g28088) );
  INVX0 U8360 ( .IN(n2663), .QN(n1701) );
  OA21X1 U8361 ( .IN1(n4684), .IN2(g4939), .IN3(n6358), .Q(n4683) );
  NOR2X0 U8362 ( .IN1(n4685), .IN2(n1590), .QN(n4684) );
  AO22X1 U8363 ( .IN1(n3030), .IN2(g4771), .IN3(n4693), .IN4(n1557), .Q(g28086) );
  INVX0 U8364 ( .IN(n2676), .QN(n1557) );
  OA21X1 U8365 ( .IN1(n4694), .IN2(g4771), .IN3(n6357), .Q(n4693) );
  NOR2X0 U8366 ( .IN1(n4695), .IN2(n3027), .QN(n4694) );
  AO22X1 U8367 ( .IN1(n3020), .IN2(g4894), .IN3(n4688), .IN4(n1700), .Q(g28087) );
  OA21X1 U8368 ( .IN1(n4689), .IN2(g4894), .IN3(n6355), .Q(n4688) );
  AO22X1 U8369 ( .IN1(n3057), .IN2(g4704), .IN3(n4707), .IN4(n1554), .Q(g28083) );
  OA21X1 U8370 ( .IN1(n4708), .IN2(g4704), .IN3(n6354), .Q(n4707) );
  AO22X1 U8371 ( .IN1(n3040), .IN2(g4760), .IN3(n4699), .IN4(n1556), .Q(g28085) );
  INVX0 U8372 ( .IN(n2680), .QN(n1556) );
  OA21X1 U8373 ( .IN1(n4700), .IN2(g4760), .IN3(n6358), .Q(n4699) );
  NOR2X0 U8374 ( .IN1(n4701), .IN2(n1564), .QN(n4700) );
  AO22X1 U8375 ( .IN1(n3081), .IN2(g4950), .IN3(n4678), .IN4(n1702), .Q(g28089) );
  INVX0 U8376 ( .IN(n2659), .QN(n1702) );
  OA21X1 U8377 ( .IN1(n4679), .IN2(g4950), .IN3(n6355), .Q(n4678) );
  NOR2X0 U8378 ( .IN1(n4680), .IN2(n1650), .QN(n4679) );
  AO22X1 U8379 ( .IN1(n3049), .IN2(test_so18), .IN3(n4703), .IN4(n1555), .Q(
        g28084) );
  INVX0 U8380 ( .IN(n2684), .QN(n1555) );
  OA21X1 U8381 ( .IN1(n4704), .IN2(test_so18), .IN3(n6354), .Q(n4703) );
  NOR2X0 U8382 ( .IN1(n4705), .IN2(n1562), .QN(n4704) );
  AO22X1 U8383 ( .IN1(n3072), .IN2(g4961), .IN3(n4673), .IN4(n1703), .Q(g28090) );
  INVX0 U8384 ( .IN(n2655), .QN(n1703) );
  OA21X1 U8385 ( .IN1(n4674), .IN2(g4961), .IN3(n6355), .Q(n4673) );
  NOR2X0 U8386 ( .IN1(n4675), .IN2(n3069), .QN(n4674) );
  AO22X1 U8387 ( .IN1(n1449), .IN2(g417), .IN3(n1448), .IN4(g446), .Q(g24209)
         );
  AO22X1 U8388 ( .IN1(n5173), .IN2(g4269), .IN3(n5262), .IN4(g4264), .Q(g21895) );
  AO21X1 U8389 ( .IN1(n5763), .IN2(g4258), .IN3(n6138), .Q(n5262) );
  AO22X1 U8390 ( .IN1(test_so72), .IN2(n5120), .IN3(n1443), .IN4(g174), .Q(
        g25601) );
  AO22X1 U8391 ( .IN1(g347), .IN2(n6123), .IN3(n4968), .IN4(g7540), .Q(g26891)
         );
  NOR2X0 U8392 ( .IN1(g347), .IN2(n6065), .QN(n4968) );
  AO22X1 U8393 ( .IN1(g4273), .IN2(n5170), .IN3(g4269), .IN4(n5171), .Q(g24280) );
  NAND2X0 U8394 ( .IN1(n6181), .IN2(n5172), .QN(n5171) );
  AO21X1 U8395 ( .IN1(n6199), .IN2(n5763), .IN3(n5173), .Q(n5170) );
  NAND3X0 U8396 ( .IN1(g4258), .IN2(n5764), .IN3(g4264), .QN(n5172) );
  AO22X1 U8397 ( .IN1(n6134), .IN2(g4527), .IN3(n4858), .IN4(n6294), .Q(g26964) );
  AO22X1 U8398 ( .IN1(n5752), .IN2(n4713), .IN3(g4515), .IN4(g4521), .Q(n4858)
         );
  AO22X1 U8399 ( .IN1(n4861), .IN2(n4864), .IN3(g4438), .IN4(n4865), .Q(g26955) );
  AO22X1 U8400 ( .IN1(g5142), .IN2(n4270), .IN3(test_so98), .IN4(n1434), .Q(
        g25706) );
  AO22X1 U8401 ( .IN1(g3835), .IN2(n4331), .IN3(test_so97), .IN4(n1438), .Q(
        g25682) );
  AO22X1 U8402 ( .IN1(g5835), .IN2(n4240), .IN3(g5841), .IN4(n1432), .Q(g25734) );
  AO22X1 U8403 ( .IN1(g6527), .IN2(n4209), .IN3(g6533), .IN4(n1430), .Q(g25762) );
  AO22X1 U8404 ( .IN1(g4145), .IN2(n4720), .IN3(g4112), .IN4(n1450), .Q(g28071) );
  INVX0 U8405 ( .IN(n4720), .QN(n1450) );
  AO21X1 U8406 ( .IN1(n4726), .IN2(n4725), .IN3(n6138), .Q(n4720) );
  AO22X1 U8407 ( .IN1(g3498), .IN2(n4346), .IN3(g3462), .IN4(n1439), .Q(g25670) );
  AO22X1 U8408 ( .IN1(g6541), .IN2(n4209), .IN3(g6505), .IN4(n1430), .Q(g25764) );
  AO22X1 U8409 ( .IN1(g5156), .IN2(n4270), .IN3(g5120), .IN4(n1434), .Q(g25708) );
  AO22X1 U8410 ( .IN1(g5503), .IN2(n4255), .IN3(g5467), .IN4(n1433), .Q(g25722) );
  AO22X1 U8411 ( .IN1(g174), .IN2(n5120), .IN3(g168), .IN4(n1443), .Q(g25600)
         );
  AO22X1 U8412 ( .IN1(g5489), .IN2(n4255), .IN3(g5495), .IN4(n1433), .Q(g25720) );
  AO22X1 U8413 ( .IN1(g6195), .IN2(n4225), .IN3(g6159), .IN4(n1431), .Q(g25750) );
  AO22X1 U8414 ( .IN1(g6181), .IN2(n4225), .IN3(g6187), .IN4(n1431), .Q(g25748) );
  AO22X1 U8415 ( .IN1(g3161), .IN2(n6131), .IN3(n3494), .IN4(n1527), .Q(g33022) );
  INVX0 U8416 ( .IN(n3500), .QN(n1527) );
  AO22X1 U8417 ( .IN1(g3484), .IN2(n4346), .IN3(g3490), .IN4(n1439), .Q(g25668) );
  AO22X1 U8418 ( .IN1(g6555), .IN2(n6133), .IN3(n3403), .IN4(n1840), .Q(g33068) );
  INVX0 U8419 ( .IN(n3404), .QN(n1840) );
  NOR2X0 U8420 ( .IN1(g6561), .IN2(n1283), .QN(n3403) );
  AO22X1 U8421 ( .IN1(g5170), .IN2(n6132), .IN3(n3443), .IN4(n1835), .Q(g33048) );
  INVX0 U8422 ( .IN(n3444), .QN(n1835) );
  NOR2X0 U8423 ( .IN1(g5176), .IN2(n1284), .QN(n3443) );
  AO22X1 U8424 ( .IN1(n6134), .IN2(g191), .IN3(n5129), .IN4(n6286), .Q(g25593)
         );
  OAI22X1 U8425 ( .IN1(n5130), .IN2(n5131), .IN3(n1989), .IN4(n5595), .QN(
        n5129) );
  AO22X1 U8426 ( .IN1(g843), .IN2(n4949), .IN3(n4950), .IN4(g812), .Q(g26898)
         );
  NAND2X0 U8427 ( .IN1(n6222), .IN2(n4952), .QN(n4949) );
  OA21X1 U8428 ( .IN1(n4951), .IN2(n1449), .IN3(g837), .Q(n4950) );
  NAND3X0 U8429 ( .IN1(g837), .IN2(n5733), .IN3(n4953), .QN(n4952) );
  AO22X1 U8430 ( .IN1(g504), .IN2(n5116), .IN3(g513), .IN4(n1442), .Q(g25611)
         );
  AO22X1 U8431 ( .IN1(g3863), .IN2(n6131), .IN3(n3478), .IN4(n2063), .Q(g33032) );
  INVX0 U8432 ( .IN(n3479), .QN(n2063) );
  NOR2X0 U8433 ( .IN1(test_so33), .IN2(n1282), .QN(n3478) );
  AO22X1 U8434 ( .IN1(g5863), .IN2(n6132), .IN3(n3423), .IN4(n2042), .Q(g33058) );
  INVX0 U8435 ( .IN(n3424), .QN(n2042) );
  NOR2X0 U8436 ( .IN1(g5869), .IN2(n1286), .QN(n3423) );
  AO22X1 U8437 ( .IN1(g3133), .IN2(n4361), .IN3(g3139), .IN4(n1440), .Q(g25654) );
  AO22X1 U8438 ( .IN1(g3849), .IN2(n4331), .IN3(g3813), .IN4(n1438), .Q(g25684) );
  AO22X1 U8439 ( .IN1(g5517), .IN2(n6132), .IN3(n3433), .IN4(n1719), .Q(g33053) );
  INVX0 U8440 ( .IN(n3434), .QN(n1719) );
  NOR2X0 U8441 ( .IN1(g5523), .IN2(n1285), .QN(n3433) );
  AO22X1 U8442 ( .IN1(g3512), .IN2(n6131), .IN3(n3488), .IN4(n1519), .Q(g33027) );
  INVX0 U8443 ( .IN(n3489), .QN(n1519) );
  NOR2X0 U8444 ( .IN1(g3518), .IN2(n1281), .QN(n3488) );
  AO22X1 U8445 ( .IN1(g3147), .IN2(n4361), .IN3(g3111), .IN4(n1440), .Q(g25656) );
  AO22X1 U8446 ( .IN1(g5849), .IN2(n4240), .IN3(g5813), .IN4(n1432), .Q(g25736) );
  AO22X1 U8447 ( .IN1(g6209), .IN2(n6133), .IN3(n3413), .IN4(n2004), .Q(g33063) );
  INVX0 U8448 ( .IN(n3414), .QN(n2004) );
  NOR2X0 U8449 ( .IN1(g6215), .IN2(n1287), .QN(n3413) );
  AO22X1 U8450 ( .IN1(g2527), .IN2(n3129), .IN3(g2533), .IN4(n1326), .Q(g33596) );
  AO22X1 U8451 ( .IN1(g1682), .IN2(n3248), .IN3(g1687), .IN4(n1348), .Q(g33547) );
  AO22X1 U8452 ( .IN1(g1816), .IN2(n3230), .IN3(g1821), .IN4(n1357), .Q(g33555) );
  AO22X1 U8453 ( .IN1(g2102), .IN2(n3190), .IN3(g2108), .IN4(n1375), .Q(g33572) );
  AO22X1 U8454 ( .IN1(g2241), .IN2(n3169), .IN3(g2246), .IN4(n1310), .Q(g33579) );
  AO22X1 U8455 ( .IN1(g1968), .IN2(n3210), .IN3(g1974), .IN4(n1366), .Q(g33564) );
  AO22X1 U8456 ( .IN1(g2259), .IN2(n3169), .IN3(test_so62), .IN4(n1310), .Q(
        g33580) );
  AO22X1 U8457 ( .IN1(g1950), .IN2(n3210), .IN3(g1955), .IN4(n1366), .Q(g33563) );
  AO22X1 U8458 ( .IN1(g324), .IN2(n6123), .IN3(n6346), .IN4(n1540), .Q(g26883)
         );
  AO22X1 U8459 ( .IN1(g2661), .IN2(n3109), .IN3(test_so48), .IN4(n1334), .Q(
        g33604) );
  AO22X1 U8460 ( .IN1(g2643), .IN2(n3109), .IN3(g2648), .IN4(n1334), .Q(g33603) );
  AO22X1 U8461 ( .IN1(g1834), .IN2(n3230), .IN3(g1840), .IN4(n1357), .Q(g33556) );
  AO22X1 U8462 ( .IN1(g2375), .IN2(n3150), .IN3(g2380), .IN4(n1318), .Q(g33587) );
  AO22X1 U8463 ( .IN1(g2509), .IN2(n3129), .IN3(g2514), .IN4(n1326), .Q(g33595) );
  AO22X1 U8464 ( .IN1(g2393), .IN2(n3150), .IN3(g2399), .IN4(n1318), .Q(g33588) );
  AO22X1 U8465 ( .IN1(g1700), .IN2(n3248), .IN3(test_so15), .IN4(n1348), .Q(
        g33548) );
  AO22X1 U8466 ( .IN1(n5981), .IN2(n5982), .IN3(n5983), .IN4(n5984), .Q(n3935)
         );
  XNOR2X1 U8467 ( .IN1(n3939), .IN2(g24181), .Q(n5982) );
  XNOR2X1 U8468 ( .IN1(n3938), .IN2(g24176), .Q(n5984) );
  AO22X1 U8469 ( .IN1(g1266), .IN2(g24247), .IN3(n5071), .IN4(g1249), .Q(
        g25630) );
  OAI21X1 U8470 ( .IN1(g1266), .IN2(n5655), .IN3(n6416), .QN(n5071) );
  AO22X1 U8471 ( .IN1(g4633), .IN2(n6125), .IN3(n1532), .IN4(n1298), .Q(g34259) );
  AO22X1 U8472 ( .IN1(g921), .IN2(g24231), .IN3(n5095), .IN4(g904), .Q(g25621)
         );
  OAI21X1 U8473 ( .IN1(g921), .IN2(n5654), .IN3(n6417), .QN(n5095) );
  AO22X1 U8474 ( .IN1(g2084), .IN2(n3190), .IN3(g2089), .IN4(n1375), .Q(g33571) );
  AO22X1 U8475 ( .IN1(n6135), .IN2(g1604), .IN3(n2975), .IN4(n6277), .Q(g33966) );
  OAI22X1 U8476 ( .IN1(n2956), .IN2(n2976), .IN3(n1343), .IN4(n5811), .QN(
        n2975) );
  INVX0 U8477 ( .IN(n2976), .QN(n1343) );
  NAND2X0 U8478 ( .IN1(n2972), .IN2(n5549), .QN(n2976) );
  AO22X1 U8479 ( .IN1(g4366), .IN2(n6124), .IN3(n6341), .IN4(n2406), .Q(g34882) );
  NAND2X0 U8480 ( .IN1(n2407), .IN2(n2408), .QN(n2406) );
  AO221X1 U8481 ( .IN1(n1390), .IN2(n5653), .IN3(n5298), .IN4(g4340), .IN5(
        n5348), .Q(n2408) );
  NAND3X0 U8482 ( .IN1(n2409), .IN2(n5348), .IN3(n2410), .QN(n2407) );
  AO22X1 U8483 ( .IN1(g3689), .IN2(n6272), .IN3(g3401), .IN4(n6137), .Q(g25663) );
  AO22X1 U8484 ( .IN1(g496), .IN2(n6274), .IN3(g1554), .IN4(n6137), .Q(g24258)
         );
  AO22X1 U8485 ( .IN1(g3338), .IN2(n6274), .IN3(g3050), .IN4(n6137), .Q(g25649) );
  AO22X1 U8486 ( .IN1(n6135), .IN2(g2165), .IN3(n2881), .IN4(n6290), .Q(g33994) );
  OAI22X1 U8487 ( .IN1(n2862), .IN2(n2882), .IN3(n1312), .IN4(n5812), .QN(
        n2881) );
  INVX0 U8488 ( .IN(n2882), .QN(n1312) );
  NAND3X0 U8489 ( .IN1(n1313), .IN2(n5514), .IN3(g2153), .QN(n2882) );
  AO22X1 U8490 ( .IN1(n6135), .IN2(g1874), .IN3(n2928), .IN4(n6287), .Q(g33980) );
  OAI22X1 U8491 ( .IN1(n2910), .IN2(n2929), .IN3(n1368), .IN4(n5813), .QN(
        n2928) );
  INVX0 U8492 ( .IN(n2929), .QN(n1368) );
  NAND3X0 U8493 ( .IN1(n2930), .IN2(n5503), .IN3(test_so8), .QN(n2929) );
  AO22X1 U8494 ( .IN1(n1379), .IN2(n6273), .IN3(g4473), .IN4(n2700), .Q(g34254) );
  INVX0 U8495 ( .IN(n2697), .QN(n1379) );
  OR4X1 U8496 ( .IN1(n5671), .IN2(n5382), .IN3(n6084), .IN4(test_so38), .Q(
        n2700) );
  AO22X1 U8497 ( .IN1(n6135), .IN2(g2433), .IN3(n2835), .IN4(n6291), .Q(g34008) );
  OAI22X1 U8498 ( .IN1(n2816), .IN2(n2836), .IN3(n1328), .IN4(n5814), .QN(
        n2835) );
  INVX0 U8499 ( .IN(n2836), .QN(n1328) );
  NAND3X0 U8500 ( .IN1(n1329), .IN2(n5523), .IN3(test_so79), .QN(n2836) );
  AO22X1 U8501 ( .IN1(g18095), .IN2(n6269), .IN3(test_so27), .IN4(n6136), .Q(
        g26962) );
  AO22X1 U8502 ( .IN1(g18095), .IN2(n6270), .IN3(g4558), .IN4(n6136), .Q(
        g26968) );
  AO22X1 U8503 ( .IN1(g5689), .IN2(n6273), .IN3(g5406), .IN4(n6136), .Q(g25715) );
  AO22X1 U8504 ( .IN1(g18096), .IN2(n6269), .IN3(g4561), .IN4(n6136), .Q(
        g26967) );
  AO22X1 U8505 ( .IN1(g4040), .IN2(n6271), .IN3(g3752), .IN4(n6136), .Q(g25677) );
  AO22X1 U8506 ( .IN1(g4473), .IN2(n6270), .IN3(g4459), .IN4(n6136), .Q(g26970) );
  AO22X1 U8507 ( .IN1(g18094), .IN2(n6268), .IN3(g4483), .IN4(n6136), .Q(
        g26961) );
  AO22X1 U8508 ( .IN1(g6035), .IN2(n6273), .IN3(g5752), .IN4(n6136), .Q(g25729) );
  AO22X1 U8509 ( .IN1(g6727), .IN2(n6270), .IN3(g6444), .IN4(n6136), .Q(g25757) );
  AO22X1 U8510 ( .IN1(g18096), .IN2(n6268), .IN3(g4489), .IN4(n6136), .Q(
        g26963) );
  AO22X1 U8511 ( .IN1(g18094), .IN2(n6272), .IN3(g4555), .IN4(n6137), .Q(
        g26966) );
  AO22X1 U8512 ( .IN1(test_so69), .IN2(n6271), .IN3(g6098), .IN4(n6136), .Q(
        g25743) );
  AO22X1 U8513 ( .IN1(n6135), .IN2(g2299), .IN3(n2858), .IN4(n6292), .Q(g34001) );
  OAI22X1 U8514 ( .IN1(n2839), .IN2(n2859), .IN3(n1320), .IN4(n5815), .QN(
        n2858) );
  INVX0 U8515 ( .IN(n2859), .QN(n1320) );
  NAND3X0 U8516 ( .IN1(n1321), .IN2(n5513), .IN3(g2287), .QN(n2859) );
  AO22X1 U8517 ( .IN1(n6135), .IN2(g2567), .IN3(n2811), .IN4(n6296), .Q(g34015) );
  OAI22X1 U8518 ( .IN1(n2792), .IN2(n2812), .IN3(n1336), .IN4(n5816), .QN(
        n2811) );
  INVX0 U8519 ( .IN(n2812), .QN(n1336) );
  NAND3X0 U8520 ( .IN1(n1337), .IN2(n5524), .IN3(g2555), .QN(n2812) );
  AO22X1 U8521 ( .IN1(g18098), .IN2(n6271), .IN3(g305), .IN4(n6137), .Q(g26881) );
  AO22X1 U8522 ( .IN1(g1146), .IN2(n5233), .IN3(g1152), .IN4(n1446), .Q(g24234) );
  AO22X1 U8523 ( .IN1(g1489), .IN2(n5211), .IN3(test_so12), .IN4(n1444), .Q(
        g24250) );
  AO22X1 U8524 ( .IN1(n6275), .IN2(n5214), .IN3(g1404), .IN4(n5215), .Q(g24248) );
  AO21X1 U8525 ( .IN1(n5217), .IN2(n5216), .IN3(n5401), .Q(n5214) );
  OR2X1 U8526 ( .IN1(n5216), .IN2(n6084), .Q(n5215) );
  NAND2X0 U8527 ( .IN1(g1404), .IN2(n5655), .QN(n5216) );
  AO22X1 U8528 ( .IN1(n6275), .IN2(n5236), .IN3(g1061), .IN4(n5237), .Q(g24232) );
  AO21X1 U8529 ( .IN1(n5239), .IN2(n5238), .IN3(n5392), .Q(n5236) );
  OR2X1 U8530 ( .IN1(n5238), .IN2(n6084), .Q(n5237) );
  NAND2X0 U8531 ( .IN1(g1061), .IN2(n5654), .QN(n5238) );
  AO22X1 U8532 ( .IN1(g2407), .IN2(n4093), .IN3(n1405), .IN4(test_so89), .Q(
        g30376) );
  INVX0 U8533 ( .IN(n4093), .QN(n1405) );
  NAND2X0 U8534 ( .IN1(n6183), .IN2(n4091), .QN(n4093) );
  AO22X1 U8535 ( .IN1(g2541), .IN2(n4081), .IN3(n1404), .IN4(g2547), .Q(g30381) );
  INVX0 U8536 ( .IN(n4081), .QN(n1404) );
  NAND2X0 U8537 ( .IN1(n6182), .IN2(n4079), .QN(n4081) );
  AO22X1 U8538 ( .IN1(g4125), .IN2(n6125), .IN3(n1437), .IN4(n5023), .Q(g25691) );
  NAND4X0 U8539 ( .IN1(n4726), .IN2(test_so11), .IN3(g4098), .IN4(n1843), .QN(
        n5023) );
  AO22X1 U8540 ( .IN1(g513), .IN2(n5116), .IN3(n1442), .IN4(g518), .Q(g25612)
         );
  AO22X1 U8541 ( .IN1(g278), .IN2(n6133), .IN3(n1422), .IN4(n5695), .Q(g28043)
         );
  AO22X1 U8542 ( .IN1(test_so12), .IN2(n5211), .IN3(n1444), .IN4(g1442), .Q(
        g24251) );
  AO22X1 U8543 ( .IN1(g2523), .IN2(n6129), .IN3(n6338), .IN4(n4082), .Q(g30380) );
  XNOR2X1 U8544 ( .IN1(n5420), .IN2(n1640), .Q(n4082) );
  AO22X1 U8545 ( .IN1(g376), .IN2(n6127), .IN3(n5122), .IN4(n6288), .Q(g25598)
         );
  OA21X1 U8546 ( .IN1(g385), .IN2(n2077), .IN3(n5121), .Q(n5122) );
  AO22X1 U8547 ( .IN1(g4281), .IN2(n6123), .IN3(n6346), .IN4(n5260), .Q(g21897) );
  AO22X1 U8548 ( .IN1(n6134), .IN2(test_so7), .IN3(n4508), .IN4(n6287), .Q(
        g29231) );
  OAI22X1 U8549 ( .IN1(n4509), .IN2(n4510), .IN3(n4511), .IN4(n5697), .QN(
        n4508) );
  NOR2X0 U8550 ( .IN1(n4509), .IN2(n4512), .QN(n4511) );
  NAND2X0 U8551 ( .IN1(n4496), .IN2(n4512), .QN(n4510) );
  AO22X1 U8552 ( .IN1(g5124), .IN2(n6124), .IN3(n6343), .IN4(n5009), .Q(g25705) );
  XNOR2X1 U8553 ( .IN1(n5427), .IN2(g32975), .Q(n5009) );
  AO22X1 U8554 ( .IN1(g2657), .IN2(n6129), .IN3(n6335), .IN4(n4070), .Q(g30385) );
  XNOR2X1 U8555 ( .IN1(n5418), .IN2(n1712), .Q(n4070) );
  AO22X1 U8556 ( .IN1(g4552), .IN2(n6128), .IN3(n2784), .IN4(n6280), .Q(g33617) );
  AO22X1 U8557 ( .IN1(g3817), .IN2(n6125), .IN3(n6347), .IN4(n5032), .Q(g25681) );
  XNOR2X1 U8558 ( .IN1(n5428), .IN2(n1907), .Q(n5032) );
  AO22X1 U8559 ( .IN1(g4515), .IN2(n6128), .IN3(n2779), .IN4(n6279), .Q(g33616) );
  AO22X1 U8560 ( .IN1(g3115), .IN2(n6125), .IN3(n6343), .IN4(n5042), .Q(g25653) );
  XNOR2X1 U8561 ( .IN1(n5423), .IN2(n1546), .Q(n5042) );
  AO22X1 U8562 ( .IN1(g6031), .IN2(n6127), .IN3(n6344), .IN4(n5151), .Q(g24345) );
  XNOR2X1 U8563 ( .IN1(g6035), .IN2(n5150), .Q(n5151) );
  AO22X1 U8564 ( .IN1(g1564), .IN2(n6126), .IN3(n5046), .IN4(n6293), .Q(g25638) );
  NOR2X0 U8565 ( .IN1(n5047), .IN2(n5048), .QN(n5046) );
  XNOR2X1 U8566 ( .IN1(n5049), .IN2(n5441), .Q(n5048) );
  AO22X1 U8567 ( .IN1(g2060), .IN2(n6128), .IN3(n6336), .IN4(n4427), .Q(g29246) );
  AO221X1 U8568 ( .IN1(n1859), .IN2(n4428), .IN3(n1856), .IN4(g2008), .IN5(
        n4429), .Q(n4427) );
  AO221X1 U8569 ( .IN1(n3585), .IN2(g2012), .IN3(n2228), .IN4(g2004), .IN5(
        n4430), .Q(n4428) );
  AO22X1 U8570 ( .IN1(g2079), .IN2(n3592), .IN3(n1857), .IN4(g2024), .Q(n4429)
         );
  AO22X1 U8571 ( .IN1(g5817), .IN2(n6124), .IN3(n6347), .IN4(n4999), .Q(g25733) );
  XNOR2X1 U8572 ( .IN1(n5429), .IN2(n1820), .Q(n4999) );
  AOI21X1 U8573 ( .IN1(n5985), .IN2(n5986), .IN3(g8342), .QN(n5038) );
  OR2X1 U8574 ( .IN1(g3451), .IN2(n5717), .Q(n5985) );
  AO22X1 U8575 ( .IN1(g6523), .IN2(n6133), .IN3(n6332), .IN4(n4211), .Q(g29308) );
  XNOR2X1 U8576 ( .IN1(n5659), .IN2(n4212), .Q(n4211) );
  AO22X1 U8577 ( .IN1(g2112), .IN2(n6132), .IN3(n6327), .IN4(n3187), .Q(g33574) );
  XNOR2X1 U8578 ( .IN1(g2116), .IN2(n3188), .Q(n3187) );
  AO22X1 U8579 ( .IN1(g1830), .IN2(n6131), .IN3(n6333), .IN4(n4142), .Q(g30355) );
  XNOR2X1 U8580 ( .IN1(n5665), .IN2(n1852), .Q(n4142) );
  AO22X1 U8581 ( .IN1(g2307), .IN2(n6130), .IN3(n6339), .IN4(n4098), .Q(g30373) );
  AO22X1 U8582 ( .IN1(g2327), .IN2(n4099), .IN3(n1743), .IN4(n4100), .Q(n4098)
         );
  NAND2X0 U8583 ( .IN1(g2331), .IN2(n5353), .QN(n4100) );
  AO22X1 U8584 ( .IN1(g2946), .IN2(n6123), .IN3(n6351), .IN4(n5253), .Q(g21901) );
  AO22X1 U8585 ( .IN1(g4180), .IN2(n5694), .IN3(n5254), .IN4(n5380), .Q(n5253)
         );
  NAND2X0 U8586 ( .IN1(n5694), .IN2(n5255), .QN(n5254) );
  AO22X1 U8587 ( .IN1(g370), .IN2(n6127), .IN3(n5124), .IN4(n6287), .Q(g25596)
         );
  OA21X1 U8588 ( .IN1(g376), .IN2(g358), .IN3(n5125), .Q(n5124) );
  AO22X1 U8589 ( .IN1(g4104), .IN2(n6131), .IN3(n6345), .IN4(n3939), .Q(g26939) );
  AO22X1 U8590 ( .IN1(g3689), .IN2(n6126), .IN3(n5186), .IN4(n6283), .Q(g24273) );
  NOR2X0 U8591 ( .IN1(g3698), .IN2(n5185), .QN(n5186) );
  AO22X1 U8592 ( .IN1(g5138), .IN2(n6133), .IN3(n6330), .IN4(n4271), .Q(g29284) );
  XNOR2X1 U8593 ( .IN1(n5658), .IN2(n4272), .Q(n4271) );
  AO22X1 U8594 ( .IN1(g4169), .IN2(n6125), .IN3(n5024), .IN4(g25689), .Q(
        g25690) );
  NOR2X0 U8595 ( .IN1(g4125), .IN2(n6077), .QN(n5024) );
  AO22X1 U8596 ( .IN1(g1882), .IN2(n6131), .IN3(n6330), .IN4(n4134), .Q(g30358) );
  AO22X1 U8597 ( .IN1(g1902), .IN2(n4135), .IN3(n1613), .IN4(n4136), .Q(n4134)
         );
  NAND2X0 U8598 ( .IN1(g1906), .IN2(n5354), .QN(n4136) );
  AO22X1 U8599 ( .IN1(g1559), .IN2(n6126), .IN3(n5050), .IN4(n6292), .Q(g25637) );
  NOR2X0 U8600 ( .IN1(n5047), .IN2(n5051), .QN(n5050) );
  OA21X1 U8601 ( .IN1(n5049), .IN2(n5441), .IN3(n5768), .Q(n5051) );
  AO22X1 U8602 ( .IN1(g1978), .IN2(n6134), .IN3(n6329), .IN4(n3207), .Q(g33566) );
  XNOR2X1 U8603 ( .IN1(g1982), .IN2(n3208), .Q(n3207) );
  AO22X1 U8604 ( .IN1(g1792), .IN2(n6129), .IN3(n6340), .IN4(n4449), .Q(g29242) );
  AO221X1 U8605 ( .IN1(n1855), .IN2(n4450), .IN3(n1852), .IN4(g1740), .IN5(
        n4451), .Q(n4449) );
  AO221X1 U8606 ( .IN1(n3621), .IN2(g1744), .IN3(n1952), .IN4(g1736), .IN5(
        n4452), .Q(n4450) );
  AO22X1 U8607 ( .IN1(g1811), .IN2(n3627), .IN3(n1853), .IN4(g1756), .Q(n4451)
         );
  AO22X1 U8608 ( .IN1(g5689), .IN2(n6127), .IN3(n5154), .IN4(n6285), .Q(g24342) );
  NOR2X0 U8609 ( .IN1(g5698), .IN2(n5153), .QN(n5154) );
  AO22X1 U8610 ( .IN1(g358), .IN2(n6127), .IN3(n6348), .IN4(n5123), .Q(g25597)
         );
  XOR2X1 U8611 ( .IN1(g370), .IN2(n2642), .Q(n5123) );
  AO22X1 U8612 ( .IN1(g1052), .IN2(n6128), .IN3(n4934), .IN4(n6293), .Q(g26914) );
  NOR2X0 U8613 ( .IN1(g979), .IN2(n4935), .QN(n4934) );
  XNOR2X1 U8614 ( .IN1(g1061), .IN2(n4936), .Q(n4935) );
  AO22X1 U8615 ( .IN1(g6727), .IN2(n6127), .IN3(n5139), .IN4(n6286), .Q(g24354) );
  NOR2X0 U8616 ( .IN1(g6736), .IN2(n5138), .QN(n5139) );
  AO22X1 U8617 ( .IN1(g5057), .IN2(n6130), .IN3(n4669), .IN4(n6288), .Q(g28092) );
  NOR2X0 U8618 ( .IN1(n3720), .IN2(n3719), .QN(n4669) );
  AO22X1 U8619 ( .IN1(g5069), .IN2(n6130), .IN3(n4671), .IN4(n6288), .Q(g28091) );
  NOR2X0 U8620 ( .IN1(n3722), .IN2(n3721), .QN(n4671) );
  AO22X1 U8621 ( .IN1(g1216), .IN2(n6127), .IN3(n5076), .IN4(n6291), .Q(g25628) );
  NOR2X0 U8622 ( .IN1(n5073), .IN2(n5077), .QN(n5076) );
  OA21X1 U8623 ( .IN1(n5075), .IN2(n5442), .IN3(n5767), .Q(n5077) );
  AO22X1 U8624 ( .IN1(g2619), .IN2(n6129), .IN3(n6337), .IN4(n4381), .Q(g29254) );
  AO221X1 U8625 ( .IN1(n1713), .IN2(n4382), .IN3(n1712), .IN4(g2567), .IN5(
        n4383), .Q(n4381) );
  AO221X1 U8626 ( .IN1(n3510), .IN2(g2571), .IN3(n1670), .IN4(g2563), .IN5(
        n4384), .Q(n4382) );
  AO22X1 U8627 ( .IN1(g2638), .IN2(n3516), .IN3(n1668), .IN4(g2583), .Q(n4383)
         );
  AO22X1 U8628 ( .IN1(g2735), .IN2(n6129), .IN3(n3730), .IN4(n4063), .Q(g30388) );
  XNOR2X1 U8629 ( .IN1(n5349), .IN2(n2049), .Q(n4063) );
  AO22X1 U8630 ( .IN1(g1844), .IN2(n6134), .IN3(n6341), .IN4(n3227), .Q(g33558) );
  XNOR2X1 U8631 ( .IN1(g1848), .IN2(n3228), .Q(n3227) );
  AO22X1 U8632 ( .IN1(g1657), .IN2(n6129), .IN3(n6340), .IN4(n4460), .Q(g29240) );
  AO221X1 U8633 ( .IN1(n1496), .IN2(g1620), .IN3(g1677), .IN4(n3645), .IN5(
        n4461), .Q(n4460) );
  AO22X1 U8634 ( .IN1(n1497), .IN2(g1604), .IN3(n1499), .IN4(n4462), .Q(n4461)
         );
  AO221X1 U8635 ( .IN1(n3639), .IN2(g1608), .IN3(n2218), .IN4(g1600), .IN5(
        n4463), .Q(n4462) );
  AO22X1 U8636 ( .IN1(test_so32), .IN2(n6124), .IN3(n5012), .IN4(n6296), .Q(
        g25702) );
  OA21X1 U8637 ( .IN1(n5013), .IN2(g5062), .IN3(n5690), .Q(n5012) );
  NOR2X0 U8638 ( .IN1(test_so32), .IN2(n5689), .QN(n5013) );
  AO22X1 U8639 ( .IN1(g142), .IN2(n6133), .IN3(n1411), .IN4(n4202), .Q(g30333)
         );
  XNOR2X1 U8640 ( .IN1(test_so73), .IN2(n4203), .Q(n4202) );
  AO22X1 U8641 ( .IN1(test_so31), .IN2(n6130), .IN3(n6332), .IN4(n3147), .Q(
        g33590) );
  XNOR2X1 U8642 ( .IN1(g2407), .IN2(n3148), .Q(n3147) );
  AO22X1 U8643 ( .IN1(g4284), .IN2(n6123), .IN3(n5259), .IN4(n6281), .Q(g21898) );
  XNOR2X1 U8644 ( .IN1(g9019), .IN2(n5258), .Q(n5259) );
  AO22X1 U8645 ( .IN1(g2741), .IN2(n6131), .IN3(n3730), .IN4(n3731), .Q(g31872) );
  AO221X1 U8646 ( .IN1(n2049), .IN2(n3562), .IN3(g2748), .IN4(n3506), .IN5(
        n3543), .Q(n3731) );
  AO22X1 U8647 ( .IN1(g5485), .IN2(n6133), .IN3(n6327), .IN4(n4256), .Q(g29290) );
  XNOR2X1 U8648 ( .IN1(n5660), .IN2(n4257), .Q(n4256) );
  AO22X1 U8649 ( .IN1(g4369), .IN2(n6125), .IN3(n6347), .IN4(n2696), .Q(g34256) );
  NAND3X0 U8650 ( .IN1(n2697), .IN2(n5765), .IN3(n2698), .QN(n2696) );
  NAND2X0 U8651 ( .IN1(g4473), .IN2(n5671), .QN(n2698) );
  AO22X1 U8652 ( .IN1(g6377), .IN2(n6127), .IN3(n6349), .IN4(n5146), .Q(g24349) );
  XNOR2X1 U8653 ( .IN1(test_so69), .IN2(n5145), .Q(n5146) );
  AO22X1 U8654 ( .IN1(g6177), .IN2(n6133), .IN3(n6327), .IN4(n4226), .Q(g29302) );
  XNOR2X1 U8655 ( .IN1(n5667), .IN2(n4227), .Q(n4226) );
  AO22X1 U8656 ( .IN1(g2485), .IN2(n6129), .IN3(n6339), .IN4(n4393), .Q(g29252) );
  AO221X1 U8657 ( .IN1(n1762), .IN2(n4394), .IN3(n1640), .IN4(g2433), .IN5(
        n4395), .Q(n4393) );
  AO221X1 U8658 ( .IN1(n3529), .IN2(g2437), .IN3(n2072), .IN4(g2429), .IN5(
        n4396), .Q(n4394) );
  AO22X1 U8659 ( .IN1(g2504), .IN2(n3535), .IN3(n1641), .IN4(g2449), .Q(n4395)
         );
  AO22X1 U8660 ( .IN1(g4849), .IN2(n6128), .IN3(n2559), .IN4(n2562), .Q(g34467) );
  XNOR2X1 U8661 ( .IN1(g4854), .IN2(n2561), .Q(n2562) );
  AO22X1 U8662 ( .IN1(g1748), .IN2(n6132), .IN3(n6332), .IN4(n4146), .Q(g30353) );
  AO22X1 U8663 ( .IN1(g1768), .IN2(n4147), .IN3(n1853), .IN4(n4148), .Q(n4146)
         );
  NAND2X0 U8664 ( .IN1(g1772), .IN2(n5352), .QN(n4148) );
  AO22X1 U8665 ( .IN1(g3480), .IN2(n6131), .IN3(n6333), .IN4(n4347), .Q(g29267) );
  XNOR2X1 U8666 ( .IN1(n5668), .IN2(n4348), .Q(n4347) );
  AO22X1 U8667 ( .IN1(g2671), .IN2(n6129), .IN3(n6334), .IN4(n3106), .Q(g33606) );
  XNOR2X1 U8668 ( .IN1(g2675), .IN2(n3107), .Q(n3106) );
  AO22X1 U8669 ( .IN1(g4235), .IN2(n6126), .IN3(n6345), .IN4(n5174), .Q(g24279) );
  XNOR2X1 U8670 ( .IN1(n5175), .IN2(n5176), .Q(n5174) );
  OA22X1 U8671 ( .IN1(g8870), .IN2(n5177), .IN3(g4235), .IN4(n5726), .Q(n5176)
         );
  AO22X1 U8672 ( .IN1(g667), .IN2(n6130), .IN3(n4525), .IN4(n4530), .Q(g29225)
         );
  XNOR2X1 U8673 ( .IN1(g671), .IN2(n1538), .Q(n4530) );
  AO22X1 U8674 ( .IN1(g2098), .IN2(n6130), .IN3(n6335), .IN4(n4118), .Q(g30365) );
  XNOR2X1 U8675 ( .IN1(n5666), .IN2(n1856), .Q(n4118) );
  AO22X1 U8676 ( .IN1(g736), .IN2(n6130), .IN3(n2404), .IN4(n4521), .Q(g29228)
         );
  XOR2X1 U8677 ( .IN1(test_so60), .IN2(n4199), .Q(n4521) );
  AO22X1 U8678 ( .IN1(g5471), .IN2(n6124), .IN3(n6342), .IN4(n5004), .Q(g25719) );
  XNOR2X1 U8679 ( .IN1(n5425), .IN2(n1755), .Q(n5004) );
  AO22X1 U8680 ( .IN1(g686), .IN2(n5110), .IN3(n1442), .IN4(g667), .Q(g25615)
         );
  AO22X1 U8681 ( .IN1(g2016), .IN2(n6131), .IN3(n6331), .IN4(n4122), .Q(g30363) );
  AO22X1 U8682 ( .IN1(test_so59), .IN2(n4123), .IN3(n1857), .IN4(n4124), .Q(
        n4122) );
  NAND2X0 U8683 ( .IN1(g2040), .IN2(n5355), .QN(n4124) );
  AO22X1 U8684 ( .IN1(g4291), .IN2(n6123), .IN3(n6352), .IN4(n5258), .Q(g21899) );
  AO22X1 U8685 ( .IN1(g4643), .IN2(n6128), .IN3(n6348), .IN4(n2580), .Q(g34459) );
  NAND2X0 U8686 ( .IN1(n2581), .IN2(n2582), .QN(n2580) );
  XNOR2X1 U8687 ( .IN1(n2583), .IN2(g4340), .Q(n2581) );
  AO22X1 U8688 ( .IN1(g2841), .IN2(n6125), .IN3(n5195), .IN4(test_so9), .Q(
        g24266) );
  NOR2X0 U8689 ( .IN1(g2712), .IN2(n6078), .QN(n5195) );
  AOI21X1 U8690 ( .IN1(n5987), .IN2(n5988), .IN3(g9741), .QN(n4995) );
  OR2X1 U8691 ( .IN1(g6148), .IN2(n5718), .Q(n5987) );
  AO22X1 U8692 ( .IN1(g2269), .IN2(n6131), .IN3(n6331), .IN4(n3166), .Q(g33582) );
  XNOR2X1 U8693 ( .IN1(g2273), .IN2(n3167), .Q(n3166) );
  AO22X1 U8694 ( .IN1(g4245), .IN2(n6123), .IN3(n5261), .IN4(n6290), .Q(g21896) );
  XNOR2X1 U8695 ( .IN1(g8839), .IN2(n5260), .Q(n5261) );
  AO22X1 U8696 ( .IN1(g222), .IN2(n6127), .IN3(n6344), .IN4(n5132), .Q(g25592)
         );
  XNOR2X1 U8697 ( .IN1(g8358), .IN2(n5133), .Q(n5132) );
  NAND2X0 U8698 ( .IN1(n5130), .IN2(n1989), .QN(n5133) );
  AO22X1 U8699 ( .IN1(g1926), .IN2(n6128), .IN3(n6337), .IN4(n4438), .Q(g29244) );
  AO221X1 U8700 ( .IN1(n1770), .IN2(n4439), .IN3(n1612), .IN4(g1874), .IN5(
        n4440), .Q(n4438) );
  AO221X1 U8701 ( .IN1(n3603), .IN2(g1878), .IN3(n1661), .IN4(g1870), .IN5(
        n4441), .Q(n4439) );
  AO22X1 U8702 ( .IN1(test_so53), .IN2(n3610), .IN3(n1613), .IN4(g1890), .Q(
        n4440) );
  AO22X1 U8703 ( .IN1(g2537), .IN2(n6130), .IN3(n6329), .IN4(n3126), .Q(g33598) );
  XNOR2X1 U8704 ( .IN1(g2541), .IN2(n3127), .Q(n3126) );
  AO22X1 U8705 ( .IN1(g6509), .IN2(n6123), .IN3(n6343), .IN4(n4989), .Q(g25761) );
  XNOR2X1 U8706 ( .IN1(n5426), .IN2(n2223), .Q(n4989) );
  AO22X1 U8707 ( .IN1(g1395), .IN2(n6129), .IN3(n4909), .IN4(n6295), .Q(g26921) );
  NOR2X0 U8708 ( .IN1(test_so68), .IN2(n4910), .QN(n4909) );
  XNOR2X1 U8709 ( .IN1(g1404), .IN2(n4911), .Q(n4910) );
  AO22X1 U8710 ( .IN1(g4239), .IN2(n6124), .IN3(n5257), .IN4(n6282), .Q(g21900) );
  NOR2X0 U8711 ( .IN1(g4297), .IN2(g10122_Tj), .QN(n5257) );
  AOI21X1 U8712 ( .IN1(n5989), .IN2(n5990), .IN3(g9817), .QN(n4990) );
  OR2X1 U8713 ( .IN1(g6494), .IN2(n5719), .Q(n5989) );
  AO22X1 U8714 ( .IN1(g4462), .IN2(n6134), .IN3(n4856), .IN4(n6294), .Q(g26969) );
  NOR2X0 U8715 ( .IN1(g4473), .IN2(test_so38), .QN(n4856) );
  AO22X1 U8716 ( .IN1(g3129), .IN2(n6130), .IN3(n6334), .IN4(n4362), .Q(g29261) );
  XNOR2X1 U8717 ( .IN1(n5661), .IN2(n4363), .Q(n4362) );
  AO22X1 U8718 ( .IN1(g5037), .IN2(n6129), .IN3(n6338), .IN4(n3707), .Q(g31900) );
  NAND3X0 U8719 ( .IN1(n3708), .IN2(n1809), .IN3(n3709), .QN(n3707) );
  NAND2X0 U8720 ( .IN1(n1824), .IN2(n5605), .QN(n3709) );
  NAND4X0 U8721 ( .IN1(n3712), .IN2(g5041), .IN3(n3711), .IN4(n3710), .QN(
        n3708) );
  AO22X1 U8722 ( .IN1(n6276), .IN2(n5860), .IN3(g333), .IN4(n6136), .Q(g26890)
         );
  AO22X1 U8723 ( .IN1(g996), .IN2(n6125), .IN3(n5223), .IN4(n6282), .Q(g24240)
         );
  OA21X1 U8724 ( .IN1(n5224), .IN2(n1740), .IN3(n5225), .Q(n5223) );
  NOR3X0 U8725 ( .IN1(g13259), .IN2(g8416), .IN3(n5084), .QN(n5224) );
  OR4X1 U8726 ( .IN1(n5084), .IN2(n5226), .IN3(g13259), .IN4(g8416), .Q(n5225)
         );
  AO22X1 U8727 ( .IN1(g3680), .IN2(n6126), .IN3(n6351), .IN4(n5188), .Q(g24272) );
  XNOR2X1 U8728 ( .IN1(g3689), .IN2(n5187), .Q(n5188) );
  AO22X1 U8729 ( .IN1(g4601), .IN2(n6123), .IN3(n2591), .IN4(n2597), .Q(g34454) );
  XNOR2X1 U8730 ( .IN1(n5274), .IN2(n2590), .Q(n2597) );
  AO22X1 U8731 ( .IN1(g5685), .IN2(n6127), .IN3(n6349), .IN4(n5156), .Q(g24341) );
  XNOR2X1 U8732 ( .IN1(g5689), .IN2(n5155), .Q(n5156) );
  AO22X1 U8733 ( .IN1(g546), .IN2(n6124), .IN3(n2404), .IN4(n5249), .Q(g24211)
         );
  NAND2X0 U8734 ( .IN1(g691), .IN2(n5486), .QN(n5249) );
  AO22X1 U8735 ( .IN1(g3466), .IN2(n6125), .IN3(n6348), .IN4(n5037), .Q(g25667) );
  XNOR2X1 U8736 ( .IN1(n5424), .IN2(n1679), .Q(n5037) );
  AO22X1 U8737 ( .IN1(g2389), .IN2(n6130), .IN3(n6333), .IN4(n4094), .Q(g30375) );
  XNOR2X1 U8738 ( .IN1(n5421), .IN2(n1742), .Q(n4094) );
  AO22X1 U8739 ( .IN1(g2173), .IN2(n6130), .IN3(n6335), .IN4(n4110), .Q(g30368) );
  AO22X1 U8740 ( .IN1(g2193), .IN2(n4111), .IN3(n1861), .IN4(n4112), .Q(n4110)
         );
  NAND2X0 U8741 ( .IN1(g2197), .IN2(n5356), .QN(n4112) );
  AO22X1 U8742 ( .IN1(g6035), .IN2(n6127), .IN3(n5149), .IN4(n6285), .Q(g24346) );
  NOR2X0 U8743 ( .IN1(test_so50), .IN2(n5148), .QN(n5149) );
  AOI21X1 U8744 ( .IN1(n5991), .IN2(n5992), .IN3(g9615), .QN(n5005) );
  OR2X1 U8745 ( .IN1(g5456), .IN2(n5720), .Q(n5991) );
  AO22X1 U8746 ( .IN1(test_so91), .IN2(n6126), .IN3(n6351), .IN4(n5193), .Q(
        g24268) );
  XNOR2X1 U8747 ( .IN1(g3338), .IN2(n5192), .Q(n5193) );
  AO22X1 U8748 ( .IN1(test_so66), .IN2(n6129), .IN3(n6339), .IN4(n4074), .Q(
        g30383) );
  AO22X1 U8749 ( .IN1(test_so34), .IN2(n4075), .IN3(n1668), .IN4(n4076), .Q(
        n4074) );
  NAND2X0 U8750 ( .IN1(g2599), .IN2(n5351), .QN(n4076) );
  AOI21X1 U8751 ( .IN1(n5993), .IN2(n5994), .IN3(g8398), .QN(n5033) );
  OR2X1 U8752 ( .IN1(g3802), .IN2(n5721), .Q(n5993) );
  AO22X1 U8753 ( .IN1(g4659), .IN2(n6128), .IN3(n2569), .IN4(n2572), .Q(g34463) );
  XNOR2X1 U8754 ( .IN1(g4664), .IN2(n2571), .Q(n2572) );
  AO22X1 U8755 ( .IN1(g4818), .IN2(n6124), .IN3(n1301), .IN4(n2762), .Q(g34033) );
  XNOR2X1 U8756 ( .IN1(n5368), .IN2(n1728), .Q(n2762) );
  AO22X1 U8757 ( .IN1(g1696), .IN2(n6132), .IN3(n6328), .IN4(n4154), .Q(g30350) );
  XNOR2X1 U8758 ( .IN1(n5417), .IN2(n1497), .Q(n4154) );
  AO22X1 U8759 ( .IN1(g3352), .IN2(n6129), .IN3(n3085), .IN4(n6278), .Q(g33610) );
  NOR2X0 U8760 ( .IN1(n3086), .IN2(n3087), .QN(n3085) );
  OA221X1 U8761 ( .IN1(n3088), .IN2(n5400), .IN3(n1590), .IN4(n3089), .IN5(
        n3090), .Q(n3087) );
  AO22X1 U8762 ( .IN1(g2441), .IN2(n6130), .IN3(n6334), .IN4(n4086), .Q(g30378) );
  AO22X1 U8763 ( .IN1(g2461), .IN2(n4087), .IN3(n1641), .IN4(n4088), .Q(n4086)
         );
  NAND2X0 U8764 ( .IN1(g2465), .IN2(n5357), .QN(n4088) );
  AO22X1 U8765 ( .IN1(g4040), .IN2(n6126), .IN3(n5181), .IN4(n6284), .Q(g24277) );
  NOR2X0 U8766 ( .IN1(g4049), .IN2(n5180), .QN(n5181) );
  AO22X1 U8767 ( .IN1(test_so11), .IN2(n6133), .IN3(n1436), .IN4(n4327), .Q(
        g29275) );
  XNOR2X1 U8768 ( .IN1(n5480), .IN2(n3942), .Q(n4327) );
  AO22X1 U8769 ( .IN1(g2351), .IN2(n6129), .IN3(n6336), .IN4(n4404), .Q(g29250) );
  AO221X1 U8770 ( .IN1(n1745), .IN2(n4405), .IN3(n1742), .IN4(g2299), .IN5(
        n4406), .Q(n4404) );
  AO221X1 U8771 ( .IN1(n3547), .IN2(g2303), .IN3(n1759), .IN4(g2295), .IN5(
        n4407), .Q(n4405) );
  AO22X1 U8772 ( .IN1(g2370), .IN2(n3554), .IN3(n1743), .IN4(g2315), .Q(n4406)
         );
  AO22X1 U8773 ( .IN1(g6163), .IN2(n6124), .IN3(n6346), .IN4(n4994), .Q(g25747) );
  XNOR2X1 U8774 ( .IN1(n5430), .IN2(n1513), .Q(n4994) );
  AOI21X1 U8775 ( .IN1(n5995), .IN2(n5996), .IN3(g9680), .QN(n5000) );
  OR2X1 U8776 ( .IN1(g5802), .IN2(n5722), .Q(n5995) );
  AO22X1 U8777 ( .IN1(g4180), .IN2(n6126), .IN3(n6341), .IN4(n5175), .Q(g21891) );
  AO22X1 U8778 ( .IN1(g5112), .IN2(n6124), .IN3(n5010), .IN4(n6298), .Q(g25703) );
  OA21X1 U8779 ( .IN1(n5011), .IN2(g5022), .IN3(n5689), .Q(n5010) );
  NOR2X0 U8780 ( .IN1(g5112), .IN2(n5690), .QN(n5011) );
  AO22X1 U8781 ( .IN1(g1221), .IN2(n6127), .IN3(n5072), .IN4(n6291), .Q(g25629) );
  NOR2X0 U8782 ( .IN1(n5073), .IN2(n5074), .QN(n5072) );
  XNOR2X1 U8783 ( .IN1(n5075), .IN2(n5442), .Q(n5074) );
  AO22X1 U8784 ( .IN1(g4332), .IN2(n6128), .IN3(n2591), .IN4(n2603), .Q(g34451) );
  XNOR2X1 U8785 ( .IN1(g4584), .IN2(n2604), .Q(n2603) );
  AO22X1 U8786 ( .IN1(g479), .IN2(n6123), .IN3(n2986), .IN4(n6280), .Q(g33962)
         );
  OA21X1 U8787 ( .IN1(n2987), .IN2(n1492), .IN3(n2988), .Q(n2986) );
  OA22X1 U8788 ( .IN1(g225), .IN2(n5962), .IN3(n6018), .IN4(g232), .Q(n2987)
         );
  AO221X1 U8789 ( .IN1(g239), .IN2(n6018), .IN3(g246), .IN4(n5962), .IN5(n6016), .Q(n2988) );
  AO22X1 U8790 ( .IN1(g518), .IN2(n6123), .IN3(n4961), .IN4(n6297), .Q(g26894)
         );
  NOR2X0 U8791 ( .IN1(n4962), .IN2(n4963), .QN(n4961) );
  OA22X1 U8792 ( .IN1(n4829), .IN2(n4964), .IN3(n1888), .IN4(n5327), .Q(n4963)
         );
  NAND2X0 U8793 ( .IN1(n4828), .IN2(n5327), .QN(n4964) );
  AO22X1 U8794 ( .IN1(g4308), .IN2(n6126), .IN3(n6350), .IN4(n5168), .Q(g24282) );
  AO22X1 U8795 ( .IN1(test_so17), .IN2(n6123), .IN3(n4967), .IN4(n6297), .Q(
        g26892) );
  NOR2X0 U8796 ( .IN1(test_so17), .IN2(n4966), .QN(n4967) );
  AO22X1 U8797 ( .IN1(g4153), .IN2(n6132), .IN3(n6344), .IN4(n3938), .Q(g26940) );
  AO22X1 U8798 ( .IN1(g832), .IN2(n6123), .IN3(n4518), .IN4(n4947), .Q(g26899)
         );
  XNOR2X1 U8799 ( .IN1(n5422), .IN2(n4814), .Q(n4947) );
  AO22X1 U8800 ( .IN1(g3831), .IN2(n6131), .IN3(n6330), .IN4(n4332), .Q(g29273) );
  XNOR2X1 U8801 ( .IN1(n5662), .IN2(n4333), .Q(n4332) );
  AOI21X1 U8802 ( .IN1(n5997), .IN2(n5998), .IN3(g8277), .QN(n5043) );
  OR2X1 U8803 ( .IN1(g3100), .IN2(n5723), .Q(n5997) );
  AO22X1 U8804 ( .IN1(g301), .IN2(n6133), .IN3(n3275), .IN4(n2707), .Q(g33537)
         );
  NOR2X0 U8805 ( .IN1(n6080), .IN2(n5724), .QN(n3275) );
  AO22X1 U8806 ( .IN1(test_so69), .IN2(n6127), .IN3(n5144), .IN4(n6285), .Q(
        g24350) );
  NOR2X0 U8807 ( .IN1(g6390), .IN2(n5143), .QN(n5144) );
  AO22X1 U8808 ( .IN1(g2255), .IN2(n6130), .IN3(n6336), .IN4(n4106), .Q(g30370) );
  XNOR2X1 U8809 ( .IN1(n5419), .IN2(n1860), .Q(n4106) );
  AO22X1 U8810 ( .IN1(g3338), .IN2(n6126), .IN3(n5191), .IN4(n6283), .Q(g24269) );
  NOR2X0 U8811 ( .IN1(g3347), .IN2(n5190), .QN(n5191) );
  AO22X1 U8812 ( .IN1(g5008), .IN2(n6125), .IN3(n1305), .IN4(n2747), .Q(g34041) );
  XNOR2X1 U8813 ( .IN1(n5367), .IN2(n1609), .Q(n2747) );
  AO22X1 U8814 ( .IN1(g5831), .IN2(n6134), .IN3(n6329), .IN4(n4241), .Q(g29296) );
  XNOR2X1 U8815 ( .IN1(n5663), .IN2(n4242), .Q(n4241) );
  AO22X1 U8816 ( .IN1(g6723), .IN2(n6127), .IN3(n6349), .IN4(n5141), .Q(g24353) );
  XNOR2X1 U8817 ( .IN1(g6727), .IN2(n5140), .Q(n5141) );
  AO22X1 U8818 ( .IN1(n6134), .IN2(g1442), .IN3(n4484), .IN4(n6286), .Q(g29236) );
  OAI22X1 U8819 ( .IN1(n4485), .IN2(n4486), .IN3(n4487), .IN4(n5696), .QN(
        n4484) );
  NOR2X0 U8820 ( .IN1(n4485), .IN2(n4488), .QN(n4487) );
  NAND2X0 U8821 ( .IN1(n4472), .IN2(n4488), .QN(n4486) );
  AO22X1 U8822 ( .IN1(g1612), .IN2(n6132), .IN3(n6328), .IN4(n4158), .Q(g30348) );
  AO22X1 U8823 ( .IN1(g1632), .IN2(n4159), .IN3(n1496), .IN4(n4160), .Q(n4158)
         );
  NAND2X0 U8824 ( .IN1(g1636), .IN2(n5362), .QN(n4160) );
  AO22X1 U8825 ( .IN1(g5339), .IN2(n6126), .IN3(n6350), .IN4(n5161), .Q(g24337) );
  XNOR2X1 U8826 ( .IN1(g25219), .IN2(n5160), .Q(n5161) );
  AO22X1 U8827 ( .IN1(g1152), .IN2(n5233), .IN3(n1446), .IN4(test_so7), .Q(
        g24235) );
  AO22X1 U8828 ( .IN1(g4512), .IN2(n6133), .IN3(n6342), .IN4(n4855), .Q(g26971) );
  NAND2X0 U8829 ( .IN1(g4531), .IN2(g4581), .QN(n4855) );
  AO22X1 U8830 ( .IN1(g4584), .IN2(n6128), .IN3(n2591), .IN4(n2602), .Q(g34452) );
  XNOR2X1 U8831 ( .IN1(n5303), .IN2(n2601), .Q(n2602) );
  AO22X1 U8832 ( .IN1(g1339), .IN2(n6125), .IN3(n5201), .IN4(n6283), .Q(g24256) );
  OA21X1 U8833 ( .IN1(n5202), .IN2(n1570), .IN3(n5203), .Q(n5201) );
  NOR3X0 U8834 ( .IN1(g13272), .IN2(g8475), .IN3(n5060), .QN(n5202) );
  OR4X1 U8835 ( .IN1(n5060), .IN2(n5204), .IN3(g13272), .IN4(g8475), .Q(n5203)
         );
  AO22X1 U8836 ( .IN1(g1964), .IN2(n6131), .IN3(n6338), .IN4(n4130), .Q(g30360) );
  XNOR2X1 U8837 ( .IN1(n5664), .IN2(n1612), .Q(n4130) );
  AO22X1 U8838 ( .IN1(g2217), .IN2(n6128), .IN3(n6340), .IN4(n4416), .Q(g29248) );
  AO221X1 U8839 ( .IN1(n1863), .IN2(n4417), .IN3(n1860), .IN4(g2165), .IN5(
        n4418), .Q(n4416) );
  AO221X1 U8840 ( .IN1(n3566), .IN2(g2169), .IN3(n2131), .IN4(g2161), .IN5(
        n4419), .Q(n4417) );
  AO22X1 U8841 ( .IN1(g2236), .IN2(n3573), .IN3(n1861), .IN4(g2181), .Q(n4418)
         );
  AO22X1 U8842 ( .IN1(g1710), .IN2(n6134), .IN3(n6331), .IN4(n3245), .Q(g33550) );
  XNOR2X1 U8843 ( .IN1(g1714), .IN2(n3246), .Q(n3245) );
  AO22X1 U8844 ( .IN1(g4031), .IN2(n6128), .IN3(n6350), .IN4(n5183), .Q(g24276) );
  XNOR2X1 U8845 ( .IN1(g4040), .IN2(n5182), .Q(n5183) );
  AO22X1 U8846 ( .IN1(n6135), .IN2(g1959), .IN3(n4131), .IN4(n6278), .Q(g30359) );
  OAI22X1 U8847 ( .IN1(n4132), .IN2(n4133), .IN3(n1660), .IN4(n5315), .QN(
        n4131) );
  XNOR2X1 U8848 ( .IN1(g1955), .IN2(g1959), .Q(n4132) );
  INVX0 U8849 ( .IN(n4133), .QN(n1660) );
  AO22X1 U8850 ( .IN1(n6135), .IN2(g1825), .IN3(n4143), .IN4(n6279), .Q(g30354) );
  OAI22X1 U8851 ( .IN1(n4144), .IN2(n4145), .IN3(n1854), .IN4(n5413), .QN(
        n4143) );
  XNOR2X1 U8852 ( .IN1(g1821), .IN2(g1825), .Q(n4144) );
  INVX0 U8853 ( .IN(n4145), .QN(n1854) );
  AO22X1 U8854 ( .IN1(n6134), .IN2(test_so78), .IN3(n4119), .IN4(n6277), .Q(
        g30364) );
  OAI22X1 U8855 ( .IN1(n4120), .IN2(n4121), .IN3(n1858), .IN4(n5280), .QN(
        n4119) );
  XNOR2X1 U8856 ( .IN1(g2089), .IN2(test_so78), .Q(n4120) );
  INVX0 U8857 ( .IN(n4121), .QN(n1858) );
  AO22X1 U8858 ( .IN1(n6135), .IN2(g2384), .IN3(n4095), .IN4(n6276), .Q(g30374) );
  OAI22X1 U8859 ( .IN1(n4096), .IN2(n4097), .IN3(n1744), .IN4(n5631), .QN(
        n4095) );
  XNOR2X1 U8860 ( .IN1(g2380), .IN2(g2384), .Q(n4096) );
  INVX0 U8861 ( .IN(n4097), .QN(n1744) );
  AO22X1 U8862 ( .IN1(n6135), .IN2(g2518), .IN3(n4083), .IN4(n6277), .Q(g30379) );
  OAI22X1 U8863 ( .IN1(n4084), .IN2(n4085), .IN3(n1761), .IN4(n5281), .QN(
        n4083) );
  XNOR2X1 U8864 ( .IN1(g2514), .IN2(g2518), .Q(n4084) );
  INVX0 U8865 ( .IN(n4085), .QN(n1761) );
  AO22X1 U8866 ( .IN1(n6134), .IN2(g1691), .IN3(n4155), .IN4(n6279), .Q(g30349) );
  OAI22X1 U8867 ( .IN1(n4156), .IN2(n4157), .IN3(n1498), .IN4(n5628), .QN(
        n4155) );
  XNOR2X1 U8868 ( .IN1(g1687), .IN2(g1691), .Q(n4156) );
  INVX0 U8869 ( .IN(n4157), .QN(n1498) );
  AO22X1 U8870 ( .IN1(n6135), .IN2(g2250), .IN3(n4107), .IN4(n6281), .Q(g30369) );
  OAI22X1 U8871 ( .IN1(n4108), .IN2(n4109), .IN3(n1862), .IN4(n5414), .QN(
        n4107) );
  XNOR2X1 U8872 ( .IN1(g2246), .IN2(g2250), .Q(n4108) );
  INVX0 U8873 ( .IN(n4109), .QN(n1862) );
  AO22X1 U8874 ( .IN1(n6135), .IN2(g2652), .IN3(n4071), .IN4(n6278), .Q(g30384) );
  OAI22X1 U8875 ( .IN1(n4072), .IN2(n4073), .IN3(n1669), .IN4(n5316), .QN(
        n4071) );
  XNOR2X1 U8876 ( .IN1(g2648), .IN2(g2652), .Q(n4072) );
  INVX0 U8877 ( .IN(n4073), .QN(n1669) );
  AO22X1 U8878 ( .IN1(g460), .IN2(n5120), .IN3(n1443), .IN4(g452), .Q(g25604)
         );
  AO22X1 U8879 ( .IN1(g1484), .IN2(n5054), .IN3(n5055), .IN4(n6292), .Q(g25635) );
  NOR2X0 U8880 ( .IN1(g1484), .IN2(n5483), .QN(n5055) );
  NAND4X0 U8881 ( .IN1(n6196), .IN2(n5056), .IN3(n5057), .IN4(n5058), .QN(
        n5054) );
  NAND2X0 U8882 ( .IN1(g1300), .IN2(n4899), .QN(n5057) );
  AO22X1 U8883 ( .IN1(g1454), .IN2(n4904), .IN3(n4905), .IN4(n6295), .Q(g26922) );
  NOR2X0 U8884 ( .IN1(g1454), .IN2(n5343), .QN(n4905) );
  NAND4X0 U8885 ( .IN1(n6198), .IN2(n4906), .IN3(n4907), .IN4(n4908), .QN(
        n4904) );
  NAND2X0 U8886 ( .IN1(g1448), .IN2(n4899), .QN(n4907) );
  AO22X1 U8887 ( .IN1(test_so90), .IN2(n4929), .IN3(n4930), .IN4(n6296), .Q(
        g26915) );
  NOR2X0 U8888 ( .IN1(test_so90), .IN2(n5478), .QN(n4930) );
  NAND4X0 U8889 ( .IN1(n6197), .IN2(n4931), .IN3(n4932), .IN4(n4933), .QN(
        n4929) );
  NAND2X0 U8890 ( .IN1(g1105), .IN2(n4924), .QN(n4932) );
  AO22X1 U8891 ( .IN1(g817), .IN2(n5097), .IN3(n5098), .IN4(g832), .Q(g25618)
         );
  NAND2X0 U8892 ( .IN1(n6187), .IN2(n5100), .QN(n5097) );
  NOR2X0 U8893 ( .IN1(n4520), .IN2(n5099), .QN(n5098) );
  OR3X1 U8894 ( .IN1(n4520), .IN2(g832), .IN3(n2076), .Q(n5100) );
  AO22X1 U8895 ( .IN1(g645), .IN2(n1421), .IN3(n4816), .IN4(g446), .Q(g28046)
         );
  AO22X1 U8896 ( .IN1(g732), .IN2(n4954), .IN3(n1428), .IN4(g753), .Q(g26897)
         );
  INVX0 U8897 ( .IN(n4954), .QN(n1428) );
  NAND2X0 U8898 ( .IN1(n6230), .IN2(n4955), .QN(n4954) );
  AO22X1 U8899 ( .IN1(g1312), .IN2(n5064), .IN3(n4914), .IN4(n5065), .Q(g25632) );
  AO21X1 U8900 ( .IN1(n4800), .IN2(n5066), .IN3(n1837), .Q(n5065) );
  NAND2X0 U8901 ( .IN1(n6201), .IN2(n5063), .QN(n5064) );
  AO22X1 U8902 ( .IN1(test_so20), .IN2(n5088), .IN3(n4939), .IN4(n5089), .Q(
        g25623) );
  AO21X1 U8903 ( .IN1(n4807), .IN2(n5090), .IN3(n1927), .Q(n5089) );
  NAND2X0 U8904 ( .IN1(n6200), .IN2(n5087), .QN(n5088) );
  AO22X1 U8905 ( .IN1(g650), .IN2(n4815), .IN3(n1421), .IN4(g655), .Q(g28050)
         );
  AO22X1 U8906 ( .IN1(g645), .IN2(n4815), .IN3(n1421), .IN4(g681), .Q(g28047)
         );
  AO22X1 U8907 ( .IN1(g655), .IN2(n4815), .IN3(n1421), .IN4(g718), .Q(g28051)
         );
  AO22X1 U8908 ( .IN1(n6134), .IN2(g446), .IN3(n2640), .IN4(n6290), .Q(g34440)
         );
  OAI22X1 U8909 ( .IN1(n2641), .IN2(n5682), .IN3(n5431), .IN4(n5305), .QN(
        n2640) );
  OA21X1 U8910 ( .IN1(n2642), .IN2(n2643), .IN3(g896), .Q(n2641) );
  NOR3X0 U8911 ( .IN1(n2644), .IN2(g703), .IN3(n2645), .QN(n2643) );
  AO22X1 U8912 ( .IN1(g661), .IN2(n4815), .IN3(n1421), .IN4(g728), .Q(g28054)
         );
  AO22X1 U8913 ( .IN1(g718), .IN2(n4815), .IN3(n1421), .IN4(g661), .Q(g28052)
         );
  AO221X1 U8914 ( .IN1(g2357), .IN2(n3098), .IN3(test_so21), .IN4(n6086), 
        .IN5(n3544), .Q(g33010) );
  OAI21X1 U8915 ( .IN1(n3545), .IN2(n6139), .IN3(n3546), .QN(n3544) );
  OA22X1 U8916 ( .IN1(n3551), .IN2(n3552), .IN3(n3553), .IN4(n5276), .Q(n3545)
         );
  NAND4X0 U8917 ( .IN1(n1745), .IN2(n3547), .IN3(n3548), .IN4(n1288), .QN(
        n3546) );
  AO221X1 U8918 ( .IN1(g2472), .IN2(n3098), .IN3(test_so79), .IN4(n6088), 
        .IN5(n3119), .Q(g33599) );
  OAI21X1 U8919 ( .IN1(n3120), .IN2(n6140), .IN3(n3121), .QN(n3119) );
  OA22X1 U8920 ( .IN1(n1295), .IN2(n3124), .IN3(n3125), .IN4(n5619), .Q(n3120)
         );
  NAND4X0 U8921 ( .IN1(n3122), .IN2(n2720), .IN3(n1288), .IN4(n3123), .QN(
        n3121) );
  AO221X1 U8922 ( .IN1(g2066), .IN2(n3098), .IN3(g2051), .IN4(n6085), .IN5(
        n3582), .Q(g33002) );
  OAI21X1 U8923 ( .IN1(n3583), .IN2(n6140), .IN3(n3584), .QN(n3582) );
  OA22X1 U8924 ( .IN1(n3589), .IN2(n3590), .IN3(n3591), .IN4(n5832), .Q(n3583)
         );
  NAND4X0 U8925 ( .IN1(n1859), .IN2(n3585), .IN3(n3586), .IN4(n1288), .QN(
        n3584) );
  AO221X1 U8926 ( .IN1(test_so75), .IN2(n3098), .IN3(g1592), .IN4(n6087), 
        .IN5(n3237), .Q(g33551) );
  OAI21X1 U8927 ( .IN1(n3238), .IN2(n6139), .IN3(n3239), .QN(n3237) );
  OA22X1 U8928 ( .IN1(n3242), .IN2(n3243), .IN3(n3244), .IN4(n5621), .Q(n3238)
         );
  NAND4X0 U8929 ( .IN1(n1474), .IN2(n3240), .IN3(g31862), .IN4(n3241), .QN(
        n3239) );
  AO221X1 U8930 ( .IN1(g1932), .IN2(n3098), .IN3(g1917), .IN4(n6085), .IN5(
        n3600), .Q(g32998) );
  OAI21X1 U8931 ( .IN1(n3601), .IN2(n6139), .IN3(n3602), .QN(n3600) );
  OA22X1 U8932 ( .IN1(n3607), .IN2(n3608), .IN3(n3609), .IN4(n5829), .Q(n3601)
         );
  NAND4X0 U8933 ( .IN1(n1770), .IN2(n3603), .IN3(n3604), .IN4(n1288), .QN(
        n3602) );
  AO221X1 U8934 ( .IN1(g2491), .IN2(n3098), .IN3(g2476), .IN4(n6086), .IN5(
        n3526), .Q(g33014) );
  OAI21X1 U8935 ( .IN1(n3527), .IN2(n6139), .IN3(n3528), .QN(n3526) );
  OA22X1 U8936 ( .IN1(n3532), .IN2(n3533), .IN3(n3534), .IN4(n5405), .Q(n3527)
         );
  NAND4X0 U8937 ( .IN1(n1762), .IN2(n3529), .IN3(n3530), .IN4(n1288), .QN(
        n3528) );
  AO221X1 U8938 ( .IN1(g1913), .IN2(n3098), .IN3(test_so8), .IN4(n6088), .IN5(
        n3198), .Q(g33567) );
  OAI21X1 U8939 ( .IN1(n3199), .IN2(n6139), .IN3(n3200), .QN(n3198) );
  OA22X1 U8940 ( .IN1(n3203), .IN2(n3204), .IN3(n3205), .IN4(n5828), .Q(n3199)
         );
  NAND4X0 U8941 ( .IN1(n3201), .IN2(n1478), .IN3(n1288), .IN4(n3202), .QN(
        n3200) );
  AO221X1 U8942 ( .IN1(g2338), .IN2(n3098), .IN3(g2287), .IN4(n6087), .IN5(
        n3138), .Q(g33591) );
  OAI21X1 U8943 ( .IN1(n3139), .IN2(n6139), .IN3(n3140), .QN(n3138) );
  OA22X1 U8944 ( .IN1(n3143), .IN2(n3144), .IN3(n3145), .IN4(n5310), .Q(n3139)
         );
  NAND4X0 U8945 ( .IN1(n3141), .IN2(n2721), .IN3(n1288), .IN4(n3142), .QN(
        n3140) );
  AO221X1 U8946 ( .IN1(g2204), .IN2(n3098), .IN3(g2153), .IN4(n6088), .IN5(
        n3157), .Q(g33583) );
  OAI21X1 U8947 ( .IN1(n3158), .IN2(n6139), .IN3(n3159), .QN(n3157) );
  OA22X1 U8948 ( .IN1(n3162), .IN2(n3163), .IN3(n3164), .IN4(n5620), .Q(n3158)
         );
  NAND4X0 U8949 ( .IN1(n3160), .IN2(n2722), .IN3(n1288), .IN4(n3161), .QN(
        n3159) );
  AO221X1 U8950 ( .IN1(test_so40), .IN2(n3098), .IN3(g2610), .IN4(n6087), 
        .IN5(n3507), .Q(g33018) );
  OAI21X1 U8951 ( .IN1(n3508), .IN2(n6139), .IN3(n3509), .QN(n3507) );
  OA22X1 U8952 ( .IN1(n3513), .IN2(n3514), .IN3(n3515), .IN4(n5277), .Q(n3508)
         );
  NAND4X0 U8953 ( .IN1(n1713), .IN2(n3510), .IN3(n3511), .IN4(n1288), .QN(
        n3509) );
  AO221X1 U8954 ( .IN1(g1779), .IN2(n3098), .IN3(g1728), .IN4(n6088), .IN5(
        n3218), .Q(g33559) );
  OAI21X1 U8955 ( .IN1(n3219), .IN2(n6139), .IN3(n3220), .QN(n3218) );
  OA22X1 U8956 ( .IN1(n3223), .IN2(n3224), .IN3(n3225), .IN4(n5830), .Q(n3219)
         );
  NAND4X0 U8957 ( .IN1(n3221), .IN2(n1476), .IN3(n1288), .IN4(n3222), .QN(
        n3220) );
  AO221X1 U8958 ( .IN1(g2047), .IN2(n3098), .IN3(g1996), .IN4(n6088), .IN5(
        n3178), .Q(g33575) );
  OAI21X1 U8959 ( .IN1(n3179), .IN2(n6139), .IN3(n3180), .QN(n3178) );
  OA22X1 U8960 ( .IN1(n3183), .IN2(n3184), .IN3(n3185), .IN4(n5831), .Q(n3179)
         );
  NAND4X0 U8961 ( .IN1(n3181), .IN2(n1480), .IN3(n1288), .IN4(n3182), .QN(
        n3180) );
  AO221X1 U8962 ( .IN1(g2223), .IN2(n3098), .IN3(g2208), .IN4(n6085), .IN5(
        n3563), .Q(g33006) );
  OAI21X1 U8963 ( .IN1(n3564), .IN2(n6139), .IN3(n3565), .QN(n3563) );
  OA22X1 U8964 ( .IN1(n3570), .IN2(n3571), .IN3(n3572), .IN4(n5406), .Q(n3564)
         );
  NAND4X0 U8965 ( .IN1(n1863), .IN2(n3566), .IN3(n3567), .IN4(n1288), .QN(
        n3565) );
  AO221X1 U8966 ( .IN1(g1664), .IN2(n3098), .IN3(test_so94), .IN4(n6084), 
        .IN5(n3636), .Q(g32990) );
  OAI21X1 U8967 ( .IN1(n3637), .IN2(n6139), .IN3(n3638), .QN(n3636) );
  OA22X1 U8968 ( .IN1(n3642), .IN2(n3643), .IN3(n3644), .IN4(n5407), .Q(n3637)
         );
  NAND4X0 U8969 ( .IN1(n1499), .IN2(n3639), .IN3(n3640), .IN4(n1288), .QN(
        n3638) );
  AO221X1 U8970 ( .IN1(g1798), .IN2(n3098), .IN3(g1783), .IN4(n6085), .IN5(
        n3618), .Q(g32994) );
  OAI21X1 U8971 ( .IN1(n3619), .IN2(n6139), .IN3(n3620), .QN(n3618) );
  OA22X1 U8972 ( .IN1(n3624), .IN2(n3625), .IN3(n3626), .IN4(n5833), .Q(n3619)
         );
  NAND4X0 U8973 ( .IN1(n1855), .IN2(n3621), .IN3(n3622), .IN4(n1288), .QN(
        n3620) );
  ISOLANDX1 U8974 ( .D(n3362), .ISO(test_so25), .Q(n2552) );
  ISOLANDX1 U8975 ( .D(n3174), .ISO(g528), .Q(n3195) );
  AO21X1 U8976 ( .IN1(n6200), .IN2(n5823), .IN3(g21893), .Q(n5173) );
  NAND4X0 U8977 ( .IN1(n1399), .IN2(g5046), .IN3(n3705), .IN4(n1809), .QN(
        n3704) );
  AO22X1 U8978 ( .IN1(g6565), .IN2(n6133), .IN3(n3398), .IN4(n3399), .Q(g33070) );
  AO221X1 U8979 ( .IN1(n2222), .IN2(n6147), .IN3(g25756), .IN4(n5646), .IN5(
        n3400), .Q(n3398) );
  AO22X1 U8980 ( .IN1(g6219), .IN2(n6133), .IN3(n3408), .IN4(n3409), .Q(g33065) );
  AO221X1 U8981 ( .IN1(n1511), .IN2(n6158), .IN3(g25742), .IN4(n5651), .IN5(
        n3410), .Q(n3408) );
  AO22X1 U8982 ( .IN1(g5180), .IN2(n6132), .IN3(n3438), .IN4(n3439), .Q(g33050) );
  AO221X1 U8983 ( .IN1(n1578), .IN2(n6160), .IN3(g25700), .IN4(n5650), .IN5(
        n3440), .Q(n3438) );
  AO22X1 U8984 ( .IN1(g3873), .IN2(n6131), .IN3(n3473), .IN4(n3474), .Q(g33034) );
  AO221X1 U8985 ( .IN1(n1905), .IN2(n6148), .IN3(g25676), .IN4(n5648), .IN5(
        n3475), .Q(n3473) );
  AO22X1 U8986 ( .IN1(g5527), .IN2(n6132), .IN3(n3428), .IN4(n3429), .Q(g33055) );
  AO221X1 U8987 ( .IN1(n1967), .IN2(n6153), .IN3(g25714), .IN4(n5647), .IN5(
        n3430), .Q(n3428) );
  AO22X1 U8988 ( .IN1(g5873), .IN2(n6133), .IN3(n3418), .IN4(n3419), .Q(g33060) );
  AO221X1 U8989 ( .IN1(n1818), .IN2(n6155), .IN3(g25728), .IN4(n5649), .IN5(
        n3420), .Q(n3418) );
  AO22X1 U8990 ( .IN1(g3522), .IN2(n6131), .IN3(n3483), .IN4(n3484), .Q(g33029) );
  AO221X1 U8991 ( .IN1(n1678), .IN2(n6154), .IN3(g25662), .IN4(n5645), .IN5(
        n3485), .Q(n3483) );
  AO221X1 U8992 ( .IN1(n4972), .IN2(g324), .IN3(g336), .IN4(n6088), .IN5(n4973), .Q(g26887) );
  NOR2X0 U8993 ( .IN1(g311), .IN2(n6065), .QN(n4972) );
  AO221X1 U8994 ( .IN1(n1877), .IN2(g24174), .IN3(g4507), .IN4(n3934), .IN5(
        n6084), .Q(g30458) );
  INVX0 U8995 ( .IN(n3934), .QN(n1877) );
  NAND2X0 U8996 ( .IN1(g4473), .IN2(n5765), .QN(n3934) );
  AO221X1 U8997 ( .IN1(n3098), .IN2(g2606), .IN3(g2555), .IN4(n6088), .IN5(
        n3099), .Q(g33607) );
  OAI21X1 U8998 ( .IN1(n3100), .IN2(n6140), .IN3(n3101), .QN(n3099) );
  OA22X1 U8999 ( .IN1(n1296), .IN2(n3104), .IN3(n3105), .IN4(n5311), .Q(n3100)
         );
  NAND4X0 U9000 ( .IN1(n3102), .IN2(n1288), .IN3(n2719), .IN4(n3103), .QN(
        n3101) );
  AO221X1 U9001 ( .IN1(n1402), .IN2(n2416), .IN3(test_so93), .IN4(n6028), 
        .IN5(n1401), .Q(g33044) );
  INVX0 U9002 ( .IN(n3453), .QN(n1401) );
  AO221X1 U9003 ( .IN1(n1402), .IN2(n2416), .IN3(g4504), .IN4(n6028), .IN5(
        n1400), .Q(g33040) );
  INVX0 U9004 ( .IN(n3462), .QN(n1400) );
  AO221X1 U9005 ( .IN1(g311), .IN2(n6149), .IN3(g316), .IN4(n6088), .IN5(n4973), .Q(g26882) );
  AO221X1 U9006 ( .IN1(n1810), .IN2(n6156), .IN3(g5041), .IN4(n6085), .IN5(
        n3702), .Q(g31901) );
  INVX0 U9007 ( .IN(n3698), .QN(n1810) );
  NAND2X0 U9008 ( .IN1(n3703), .IN2(n3704), .QN(n3702) );
  NAND2X0 U9009 ( .IN1(n1823), .IN2(n5578), .QN(n3703) );
  AO221X1 U9010 ( .IN1(n1449), .IN2(test_so87), .IN3(g681), .IN4(n6087), .IN5(
        n4816), .Q(g28053) );
  AO221X1 U9011 ( .IN1(n3688), .IN2(n6163), .IN3(g5029), .IN4(n6085), .IN5(
        n3689), .Q(g31904) );
  NAND2X0 U9012 ( .IN1(n3690), .IN2(n3691), .QN(n3689) );
  OR2X1 U9013 ( .IN1(n3692), .IN2(g5033), .Q(n3690) );
  NAND4X0 U9014 ( .IN1(n1399), .IN2(g5033), .IN3(n3692), .IN4(n3693), .QN(
        n3691) );
  AO221X1 U9015 ( .IN1(n6159), .IN2(n4827), .IN3(g528), .IN4(n6087), .IN5(
        n1441), .Q(g28044) );
  XNOR2X1 U9016 ( .IN1(g482), .IN2(n4542), .Q(n4827) );
  AO221X1 U9017 ( .IN1(g2197), .IN2(n2863), .IN3(g2204), .IN4(n6088), .IN5(
        n3171), .Q(g33577) );
  NOR4X0 U9018 ( .IN1(n1293), .IN2(n2870), .IN3(n6115), .IN4(n5356), .QN(n3171) );
  AO221X1 U9019 ( .IN1(g2331), .IN2(n2840), .IN3(g2338), .IN4(n6088), .IN5(
        n3152), .Q(g33585) );
  NOR4X0 U9020 ( .IN1(n1294), .IN2(n2847), .IN3(n6116), .IN4(n5353), .QN(n3152) );
  AO221X1 U9021 ( .IN1(n6150), .IN2(n4887), .IN3(g4141), .IN4(n6088), .IN5(
        n1437), .Q(g26938) );
  XOR2X1 U9022 ( .IN1(g4082), .IN2(n4729), .Q(n4887) );
  AO221X1 U9023 ( .IN1(g1906), .IN2(n2911), .IN3(g1913), .IN4(n6087), .IN5(
        n3212), .Q(g33561) );
  NOR4X0 U9024 ( .IN1(n1291), .IN2(n1365), .IN3(n6115), .IN4(n5354), .QN(n3212) );
  AO221X1 U9025 ( .IN1(g2040), .IN2(n2887), .IN3(g2047), .IN4(n6087), .IN5(
        n3192), .Q(g33569) );
  NOR4X0 U9026 ( .IN1(n1292), .IN2(n1374), .IN3(n6115), .IN4(n5355), .QN(n3192) );
  AO221X1 U9027 ( .IN1(g703), .IN2(n5245), .IN3(g847), .IN4(n6086), .IN5(n5246), .Q(g24214) );
  NOR4X0 U9028 ( .IN1(n5422), .IN2(n5247), .IN3(n5826), .IN4(n5102), .QN(n5246) );
  NAND2X0 U9029 ( .IN1(n4545), .IN2(n5248), .QN(n5245) );
  AO221X1 U9030 ( .IN1(n1645), .IN2(n5715), .IN3(g4098), .IN4(n6087), .IN5(
        n3468), .Q(g33035) );
  NAND2X0 U9031 ( .IN1(n3469), .IN2(n3470), .QN(n3468) );
  NAND3X0 U9032 ( .IN1(n6417), .IN2(n3471), .IN3(g4108), .QN(n3469) );
  AO221X1 U9033 ( .IN1(n3452), .IN2(n6161), .IN3(g5046), .IN4(n6085), .IN5(
        n3694), .Q(g31903) );
  NAND2X0 U9034 ( .IN1(n3695), .IN2(n3696), .QN(n3694) );
  NAND2X0 U9035 ( .IN1(n1822), .IN2(n5607), .QN(n3695) );
  NAND4X0 U9036 ( .IN1(n1399), .IN2(g5052), .IN3(n3697), .IN4(n3698), .QN(
        n3696) );
  AO221X1 U9037 ( .IN1(g1772), .IN2(n2934), .IN3(g1779), .IN4(n6087), .IN5(
        n3232), .Q(g33553) );
  NOR4X0 U9038 ( .IN1(n1290), .IN2(n1356), .IN3(n6115), .IN4(n5352), .QN(n3232) );
  AO221X1 U9039 ( .IN1(g2599), .IN2(n2793), .IN3(g2606), .IN4(n6088), .IN5(
        n3112), .Q(g33601) );
  NOR4X0 U9040 ( .IN1(n3111), .IN2(n2800), .IN3(n6116), .IN4(n5351), .QN(n3112) );
  AO221X1 U9041 ( .IN1(n6151), .IN2(n3728), .IN3(g4093), .IN4(n6086), .IN5(
        n1437), .Q(g31894) );
  XNOR2X1 U9042 ( .IN1(n5350), .IN2(n3472), .Q(n3728) );
  AO221X1 U9043 ( .IN1(g2465), .IN2(n2817), .IN3(g2472), .IN4(n6087), .IN5(
        n3132), .Q(g33593) );
  NOR4X0 U9044 ( .IN1(n3131), .IN2(n2824), .IN3(n6116), .IN4(n5357), .QN(n3132) );
  AO221X1 U9045 ( .IN1(n2108), .IN2(n5543), .IN3(g4082), .IN4(n6086), .IN5(
        n4727), .Q(g28070) );
  INVX0 U9046 ( .IN(n4328), .QN(n2108) );
  NAND2X0 U9047 ( .IN1(n4728), .IN2(n3470), .QN(n4727) );
  NAND3X0 U9048 ( .IN1(n6416), .IN2(n4328), .IN3(test_so11), .QN(n4728) );
  AO221X1 U9049 ( .IN1(n5232), .IN2(g1178), .IN3(g1183), .IN4(n6086), .IN5(
        n5078), .Q(g24236) );
  NOR2X0 U9050 ( .IN1(n6021), .IN2(n6077), .QN(n5232) );
  AO221X1 U9051 ( .IN1(n4538), .IN2(n5708), .IN3(g482), .IN4(n6085), .IN5(
        n4539), .Q(g29223) );
  NAND2X0 U9052 ( .IN1(n4540), .IN2(n4541), .QN(n4539) );
  OR3X1 U9053 ( .IN1(n6115), .IN2(n4538), .IN3(n5708), .Q(n4540) );
  AO21X1 U9054 ( .IN1(n2907), .IN2(n2908), .IN3(n1378), .Q(n2893) );
  NAND2X0 U9055 ( .IN1(g956), .IN2(n5286), .QN(n2908) );
  AO21X1 U9056 ( .IN1(n2907), .IN2(n2977), .IN3(n1351), .Q(n2963) );
  NAND2X0 U9057 ( .IN1(g1135), .IN2(n5286), .QN(n2977) );
  AO21X1 U9058 ( .IN1(n2907), .IN2(n2954), .IN3(n1360), .Q(n2940) );
  NAND2X0 U9059 ( .IN1(g1105), .IN2(n5286), .QN(n2954) );
  AO21X1 U9060 ( .IN1(n2907), .IN2(n2931), .IN3(n1369), .Q(n2917) );
  NAND2X0 U9061 ( .IN1(g1129), .IN2(n5286), .QN(n2931) );
  AO221X1 U9062 ( .IN1(g4072), .IN2(n6088), .IN3(n6178), .IN4(n5416), .IN5(
        n1437), .Q(g25685) );
  NAND3X0 U9063 ( .IN1(g518), .IN2(n3116), .IN3(g504), .QN(n2727) );
  NAND3X0 U9064 ( .IN1(n3116), .IN2(n5519), .IN3(g518), .QN(n2726) );
  ISOLANDX1 U9065 ( .D(g4145), .ISO(n6144), .Q(n4721) );
  NAND4X0 U9066 ( .IN1(g24162), .IN2(n5325), .IN3(n4854), .IN4(n5948), .QN(
        n3309) );
  NOR2X0 U9067 ( .IN1(g24164), .IN2(g24163), .QN(n4854) );
  OA21X1 U9068 ( .IN1(n2587), .IN2(test_so3), .IN3(n1297), .Q(n2588) );
  NAND2X0 U9069 ( .IN1(g3115), .IN2(n6148), .QN(n2473) );
  ISOLANDX1 U9070 ( .D(g2841), .ISO(n6145), .Q(n3730) );
  NAND2X0 U9071 ( .IN1(g6509), .IN2(n6177), .QN(n2474) );
  OR2X1 U9072 ( .IN1(n3344), .IN2(g1291), .Q(n3306) );
  OR2X1 U9073 ( .IN1(n3345), .IN2(g947), .Q(n3307) );
  AO21X1 U9074 ( .IN1(g385), .IN2(n6119), .IN3(n2642), .Q(g25599) );
  ISOLANDX1 U9075 ( .D(g19), .ISO(g9), .Q(n3362) );
  ISOLANDX1 U9076 ( .D(g24174), .ISO(n6144), .Q(g25694) );
  AO22X1 U9077 ( .IN1(n6275), .IN2(test_so47), .IN3(n4860), .IN4(g4434), .Q(
        g26957) );
  AO21X1 U9078 ( .IN1(g4392), .IN2(n4861), .IN3(n6137), .Q(n4860) );
  AO21X1 U9079 ( .IN1(g2984), .IN2(n1802), .IN3(n3350), .Q(n3393) );
  ISOLANDX1 U9080 ( .D(n4305), .ISO(n6144), .Q(g29277) );
  NAND3X0 U9081 ( .IN1(n4306), .IN2(n4307), .IN3(n4308), .QN(n4305) );
  OR2X1 U9082 ( .IN1(n5656), .IN2(g4826), .Q(n4307) );
  AOI222X1 U9083 ( .IN1(g4681), .IN2(g4831), .IN3(g4646), .IN4(g21245), .IN5(
        n5880), .IN6(g4674), .QN(n4308) );
  ISOLANDX1 U9084 ( .D(g4423), .ISO(n6144), .Q(g26953) );
  ISOLANDX1 U9085 ( .D(g24165), .ISO(n6144), .Q(g24212) );
  ISOLANDX1 U9086 ( .D(n4283), .ISO(n6144), .Q(g29279) );
  NAND3X0 U9087 ( .IN1(n4284), .IN2(n4285), .IN3(n4286), .QN(n4283) );
  NAND2X0 U9088 ( .IN1(g5011), .IN2(g4836), .QN(n4285) );
  OA222X1 U9089 ( .IN1(g4035), .IN2(n5283), .IN3(g3333), .IN4(n5318), .IN5(
        n5443), .IN6(n5881), .Q(n4286) );
  ISOLANDX1 U9090 ( .D(g24180), .ISO(n6145), .Q(g25688) );
  NOR4X0 U9091 ( .IN1(n5207), .IN2(g17320), .IN3(g17423), .IN4(g17404), .QN(
        g24254) );
  AO21X1 U9092 ( .IN1(n5047), .IN2(n5208), .IN3(n6137), .Q(n5207) );
  NAND3X0 U9093 ( .IN1(n4176), .IN2(n5466), .IN3(n1571), .QN(n5208) );
  AO21X1 U9094 ( .IN1(g1585), .IN2(n6121), .IN3(n1445), .Q(g24261) );
  AO21X1 U9095 ( .IN1(g4382), .IN2(n6120), .IN3(n1288), .Q(g31895) );
  AO21X1 U9096 ( .IN1(g2771), .IN2(n6119), .IN3(n4044), .Q(g30391) );
  AO21X1 U9097 ( .IN1(g2803), .IN2(n6119), .IN3(n4043), .Q(g30392) );
  ISOLANDX1 U9098 ( .D(g4681), .ISO(n2774), .Q(g34028) );
  ISOLANDX1 U9099 ( .D(n2595), .ISO(n2608), .Q(g34449) );
  XNOR2X1 U9100 ( .IN1(g4311), .IN2(n2607), .Q(n2608) );
  ISOLANDX1 U9101 ( .D(g18099), .ISO(n6144), .Q(g26880) );
  AO21X1 U9102 ( .IN1(g2831), .IN2(n6119), .IN3(n4044), .Q(g30389) );
  AO21X1 U9103 ( .IN1(g2834), .IN2(n6119), .IN3(n4043), .Q(g30390) );
  AO22X1 U9104 ( .IN1(g1811), .IN2(n4445), .IN3(n4446), .IN4(g1825), .Q(g29243) );
  OA21X1 U9105 ( .IN1(n4447), .IN2(n3627), .IN3(n6362), .Q(n4446) );
  AO21X1 U9106 ( .IN1(n1855), .IN2(n4448), .IN3(n6138), .Q(n4445) );
  ISOLANDX1 U9107 ( .D(n4448), .ISO(n1952), .Q(n4447) );
  AO22X1 U9108 ( .IN1(g2370), .IN2(n4400), .IN3(n4401), .IN4(g2384), .Q(g29251) );
  OA21X1 U9109 ( .IN1(n4402), .IN2(n3554), .IN3(n6359), .Q(n4401) );
  AO21X1 U9110 ( .IN1(n1745), .IN2(n4403), .IN3(n6138), .Q(n4400) );
  ISOLANDX1 U9111 ( .D(n4403), .ISO(n1759), .Q(n4402) );
  NOR3X0 U9112 ( .IN1(test_so85), .IN2(g8), .IN3(g6), .QN(n3396) );
  AO22X1 U9113 ( .IN1(g2079), .IN2(n4423), .IN3(n4424), .IN4(test_so78), .Q(
        g29247) );
  OA21X1 U9114 ( .IN1(n4425), .IN2(n3592), .IN3(n6358), .Q(n4424) );
  AO21X1 U9115 ( .IN1(n1859), .IN2(n4426), .IN3(n6138), .Q(n4423) );
  ISOLANDX1 U9116 ( .D(n4426), .ISO(n2228), .Q(n4425) );
  AO22X1 U9117 ( .IN1(test_so53), .IN2(n4434), .IN3(n4435), .IN4(g1959), .Q(
        g29245) );
  OA21X1 U9118 ( .IN1(n4436), .IN2(n3610), .IN3(n6357), .Q(n4435) );
  AO21X1 U9119 ( .IN1(n1770), .IN2(n4437), .IN3(n6138), .Q(n4434) );
  ISOLANDX1 U9120 ( .D(n4437), .ISO(n1661), .Q(n4436) );
  AO22X1 U9121 ( .IN1(g2504), .IN2(n4389), .IN3(n4390), .IN4(g2518), .Q(g29253) );
  OA21X1 U9122 ( .IN1(n4391), .IN2(n3535), .IN3(n6360), .Q(n4390) );
  AO21X1 U9123 ( .IN1(n1762), .IN2(n4392), .IN3(n6138), .Q(n4389) );
  ISOLANDX1 U9124 ( .D(n4392), .ISO(n2072), .Q(n4391) );
  AO22X1 U9125 ( .IN1(g2638), .IN2(n4377), .IN3(n4378), .IN4(g2652), .Q(g29255) );
  OA21X1 U9126 ( .IN1(n4379), .IN2(n3516), .IN3(n6361), .Q(n4378) );
  AO21X1 U9127 ( .IN1(n1713), .IN2(n4380), .IN3(n6138), .Q(n4377) );
  ISOLANDX1 U9128 ( .D(n4380), .ISO(n1670), .Q(n4379) );
  AO22X1 U9129 ( .IN1(g2236), .IN2(n4412), .IN3(n4413), .IN4(g2250), .Q(g29249) );
  OA21X1 U9130 ( .IN1(n4414), .IN2(n3573), .IN3(n6363), .Q(n4413) );
  AO21X1 U9131 ( .IN1(n1863), .IN2(n4415), .IN3(n6138), .Q(n4412) );
  ISOLANDX1 U9132 ( .D(n4415), .ISO(n2131), .Q(n4414) );
  AO22X1 U9133 ( .IN1(g1677), .IN2(n4456), .IN3(n4457), .IN4(g1691), .Q(g29241) );
  OA21X1 U9134 ( .IN1(n4458), .IN2(n3645), .IN3(n6356), .Q(n4457) );
  AO21X1 U9135 ( .IN1(n1499), .IN2(n4459), .IN3(n6138), .Q(n4456) );
  ISOLANDX1 U9136 ( .D(n4459), .ISO(n2218), .Q(n4458) );
  AO21X1 U9137 ( .IN1(n6201), .IN2(n4868), .IN3(n4869), .Q(g26952) );
  XOR2X1 U9138 ( .IN1(g4434), .IN2(g4401), .Q(n4868) );
  XNOR2X1 U9139 ( .IN1(g4430), .IN2(n4870), .Q(n4869) );
  NAND2X0 U9140 ( .IN1(g4388), .IN2(n6174), .QN(n4870) );
  AO21X1 U9141 ( .IN1(g1236), .IN2(n6122), .IN3(n1447), .Q(g24243) );
  AO21X1 U9142 ( .IN1(g4427), .IN2(n6120), .IN3(g26953), .Q(g26951) );
  AO21X1 U9143 ( .IN1(g1579), .IN2(n6121), .IN3(n1445), .Q(g24259) );
  AO21X1 U9144 ( .IN1(g4492), .IN2(n6120), .IN3(n2776), .Q(g34024) );
  OA221X1 U9145 ( .IN1(n2777), .IN2(n2778), .IN3(n1490), .IN4(n2779), .IN5(
        n6228), .Q(n2776) );
  AO21X1 U9146 ( .IN1(g355), .IN2(n6120), .IN3(n4965), .Q(g26893) );
  OA221X1 U9147 ( .IN1(test_so17), .IN2(g20763), .IN3(n1757), .IN4(n5825), 
        .IN5(n6230), .Q(n4965) );
  INVX0 U9148 ( .IN(n4966), .QN(n1757) );
  AO21X1 U9149 ( .IN1(g4572), .IN2(n6121), .IN3(g29279), .Q(g29278) );
  AO21X1 U9150 ( .IN1(g753), .IN2(n6122), .IN3(g24212), .Q(g24213) );
  OA21X1 U9151 ( .IN1(g1589), .IN2(n2798), .IN3(n2799), .Q(n2797) );
  OA21X1 U9152 ( .IN1(g1589), .IN2(n2845), .IN3(n2846), .Q(n2844) );
  OA21X1 U9153 ( .IN1(n6117), .IN2(n5096), .IN3(g837), .Q(g25619) );
  XOR2X1 U9154 ( .IN1(g843), .IN2(n4953), .Q(n5096) );
  OA21X1 U9155 ( .IN1(g1246), .IN2(n2892), .IN3(n2893), .Q(n2891) );
  OA21X1 U9156 ( .IN1(g1246), .IN2(n2939), .IN3(n2940), .Q(n2938) );
  NAND2X0 U9157 ( .IN1(n5218), .IN2(n5219), .QN(g24246) );
  AO21X1 U9158 ( .IN1(n5220), .IN2(n6203), .IN3(n5547), .Q(n5218) );
  NAND3X0 U9159 ( .IN1(n6416), .IN2(n5547), .IN3(g1221), .QN(n5219) );
  XNOR2X1 U9160 ( .IN1(g1087), .IN2(g1221), .Q(n5220) );
  NAND2X0 U9161 ( .IN1(n5196), .IN2(n5197), .QN(g24262) );
  AO21X1 U9162 ( .IN1(n5198), .IN2(n6204), .IN3(n5546), .Q(n5196) );
  NAND3X0 U9163 ( .IN1(n6418), .IN2(n5546), .IN3(g1564), .QN(n5197) );
  XNOR2X1 U9164 ( .IN1(g1430), .IN2(g1564), .Q(n5198) );
  NAND2X0 U9165 ( .IN1(n5819), .IN2(n4862), .QN(g26956) );
  NAND3X0 U9166 ( .IN1(n4863), .IN2(n4861), .IN3(g4430), .QN(n4862) );
  NAND2X0 U9167 ( .IN1(n2837), .IN2(n2822), .QN(n2823) );
  AO21X1 U9168 ( .IN1(g1472), .IN2(n2549), .IN3(n2814), .Q(n2837) );
  NAND2X0 U9169 ( .IN1(n2883), .IN2(n2868), .QN(n2869) );
  AO21X1 U9170 ( .IN1(g1478), .IN2(n2549), .IN3(n2814), .Q(n2883) );
  NAND2X0 U9171 ( .IN1(n2813), .IN2(n2798), .QN(n2799) );
  AO21X1 U9172 ( .IN1(g1300), .IN2(n2549), .IN3(n2814), .Q(n2813) );
  NAND2X0 U9173 ( .IN1(n2860), .IN2(n2845), .QN(n2846) );
  AO21X1 U9174 ( .IN1(g1448), .IN2(n2549), .IN3(n2814), .Q(n2860) );
  OA21X1 U9175 ( .IN1(n2710), .IN2(n6118), .IN3(g160), .Q(g33536) );
  AO21X1 U9176 ( .IN1(g1592), .IN2(n2957), .IN3(n3251), .Q(g33544) );
  NOR4X0 U9177 ( .IN1(g1668), .IN2(n1289), .IN3(n3252), .IN4(n6117), .QN(n3251) );
  OA21X1 U9178 ( .IN1(g1636), .IN2(n1347), .IN3(n5362), .Q(n3252) );
  AO21X1 U9179 ( .IN1(g2555), .IN2(n2793), .IN3(n3113), .Q(g33600) );
  NOR4X0 U9180 ( .IN1(g2629), .IN2(n3111), .IN3(n3114), .IN4(n6118), .QN(n3113) );
  OA21X1 U9181 ( .IN1(g2599), .IN2(n2800), .IN3(n5351), .Q(n3114) );
  AO21X1 U9182 ( .IN1(g1728), .IN2(n2934), .IN3(n3233), .Q(g33552) );
  NOR4X0 U9183 ( .IN1(g1802), .IN2(n1290), .IN3(n3234), .IN4(n6117), .QN(n3233) );
  OA21X1 U9184 ( .IN1(g1772), .IN2(n1356), .IN3(n5352), .Q(n3234) );
  AO21X1 U9185 ( .IN1(g2287), .IN2(n2840), .IN3(n3153), .Q(g33584) );
  NOR4X0 U9186 ( .IN1(g2361), .IN2(n1294), .IN3(n3154), .IN4(n6117), .QN(n3153) );
  OA21X1 U9187 ( .IN1(g2331), .IN2(n2847), .IN3(n5353), .Q(n3154) );
  AO21X1 U9188 ( .IN1(test_so8), .IN2(n2911), .IN3(n3213), .Q(g33560) );
  NOR4X0 U9189 ( .IN1(g1936), .IN2(n1291), .IN3(n3214), .IN4(n6117), .QN(n3213) );
  OA21X1 U9190 ( .IN1(g1906), .IN2(n1365), .IN3(n5354), .Q(n3214) );
  OAI22X1 U9191 ( .IN1(n6312), .IN2(n5683), .IN3(n2900), .IN4(n6143), .QN(
        g33989) );
  OA22X1 U9192 ( .IN1(n2886), .IN2(n2901), .IN3(n1372), .IN4(n5852), .Q(n2900)
         );
  INVX0 U9193 ( .IN(n2901), .QN(n1372) );
  OAI22X1 U9194 ( .IN1(n6315), .IN2(n5797), .IN3(n2947), .IN4(n6143), .QN(
        g33975) );
  OA22X1 U9195 ( .IN1(n2933), .IN2(n2948), .IN3(n1354), .IN4(n5853), .Q(n2947)
         );
  INVX0 U9196 ( .IN(n2948), .QN(n1354) );
  OAI22X1 U9197 ( .IN1(n6313), .IN2(n5686), .IN3(n2924), .IN4(n6142), .QN(
        g33982) );
  OA22X1 U9198 ( .IN1(n2910), .IN2(n2925), .IN3(n1363), .IN4(n5854), .Q(n2924)
         );
  INVX0 U9199 ( .IN(n2925), .QN(n1363) );
  OAI221X1 U9200 ( .IN1(n4368), .IN2(n5742), .IN3(n4363), .IN4(n2473), .IN5(
        n4369), .QN(g29258) );
  NAND4X0 U9201 ( .IN1(g3111), .IN2(n4363), .IN3(n6175), .IN4(n5742), .QN(
        n4369) );
  OA21X1 U9202 ( .IN1(g3111), .IN2(n1589), .IN3(n6366), .Q(n4368) );
  OAI221X1 U9203 ( .IN1(n5007), .IN2(n5444), .IN3(n4270), .IN4(n5883), .IN5(
        n5008), .QN(g25707) );
  NAND4X0 U9204 ( .IN1(g32975), .IN2(n6186), .IN3(n5658), .IN4(n5444), .QN(
        n5008) );
  OA21X1 U9205 ( .IN1(n3287), .IN2(n5658), .IN3(n6360), .Q(n5007) );
  OAI221X1 U9206 ( .IN1(n4277), .IN2(n5743), .IN3(n4272), .IN4(n3764), .IN5(
        n4278), .QN(g29281) );
  NAND4X0 U9207 ( .IN1(g5120), .IN2(n4272), .IN3(n6174), .IN4(n5743), .QN(
        n4278) );
  OA21X1 U9208 ( .IN1(g5120), .IN2(n1559), .IN3(n6368), .Q(n4277) );
  OAI221X1 U9209 ( .IN1(n4262), .IN2(n5744), .IN3(n4257), .IN4(n3758), .IN5(
        n4263), .QN(g29287) );
  NAND4X0 U9210 ( .IN1(g5467), .IN2(n4257), .IN3(n6169), .IN4(n5744), .QN(
        n4263) );
  OA21X1 U9211 ( .IN1(g5467), .IN2(n1561), .IN3(n6370), .Q(n4262) );
  OAI221X1 U9212 ( .IN1(n4338), .IN2(n5745), .IN3(n4333), .IN4(n2478), .IN5(
        n4339), .QN(g29270) );
  NAND4X0 U9213 ( .IN1(g3813), .IN2(n4333), .IN3(n6171), .IN4(n5745), .QN(
        n4339) );
  OA21X1 U9214 ( .IN1(g3813), .IN2(n1502), .IN3(n6366), .Q(n4338) );
  OAI221X1 U9215 ( .IN1(n4353), .IN2(n5746), .IN3(n4348), .IN4(n2475), .IN5(
        n4354), .QN(g29264) );
  NAND4X0 U9216 ( .IN1(g3462), .IN2(n4348), .IN3(n6176), .IN4(n5746), .QN(
        n4354) );
  OA21X1 U9217 ( .IN1(g3462), .IN2(n1594), .IN3(n6368), .Q(n4353) );
  OAI221X1 U9218 ( .IN1(n4987), .IN2(n5445), .IN3(n4209), .IN4(n5884), .IN5(
        n4988), .QN(g25763) );
  NAND4X0 U9219 ( .IN1(n2223), .IN2(n6190), .IN3(n5659), .IN4(n5445), .QN(
        n4988) );
  OA21X1 U9220 ( .IN1(n3295), .IN2(n5659), .IN3(n6356), .Q(n4987) );
  OAI221X1 U9221 ( .IN1(n5002), .IN2(n5446), .IN3(n4255), .IN4(n5885), .IN5(
        n5003), .QN(g25721) );
  NAND4X0 U9222 ( .IN1(n1755), .IN2(n6191), .IN3(n5660), .IN4(n5446), .QN(
        n5003) );
  OA21X1 U9223 ( .IN1(n3289), .IN2(n5660), .IN3(n6365), .Q(n5002) );
  OAI221X1 U9224 ( .IN1(n5040), .IN2(n5447), .IN3(n4361), .IN4(n5882), .IN5(
        n5041), .QN(g25655) );
  NAND4X0 U9225 ( .IN1(n1546), .IN2(n6179), .IN3(n5661), .IN4(n5447), .QN(
        n5041) );
  OA21X1 U9226 ( .IN1(n3296), .IN2(n5661), .IN3(n6363), .Q(n5040) );
  OAI22X1 U9227 ( .IN1(n2584), .IN2(n5844), .IN3(n2585), .IN4(n5309), .QN(
        g34458) );
  OA21X1 U9228 ( .IN1(g4633), .IN2(n2586), .IN3(n6364), .Q(n2585) );
  OA21X1 U9229 ( .IN1(test_so99), .IN2(n2587), .IN3(n2588), .Q(n2584) );
  OAI22X1 U9230 ( .IN1(n3497), .IN2(n5652), .IN3(n3498), .IN4(n3499), .QN(
        g33023) );
  NAND2X0 U9231 ( .IN1(g3171), .IN2(n5652), .QN(n3499) );
  OA21X1 U9232 ( .IN1(g3171), .IN2(n1280), .IN3(n6407), .Q(n3497) );
  OA22X1 U9233 ( .IN1(n5735), .IN2(n4329), .IN3(n4330), .IN4(n6047), .Q(g29274) );
  NAND2X0 U9234 ( .IN1(n4210), .IN2(n3298), .QN(n4329) );
  NOR2X0 U9235 ( .IN1(n4331), .IN2(n5735), .QN(n4330) );
  OA22X1 U9236 ( .IN1(n5736), .IN2(n4238), .IN3(n4239), .IN4(n6047), .Q(g29297) );
  NAND2X0 U9237 ( .IN1(n4210), .IN2(n3294), .QN(n4238) );
  NOR2X0 U9238 ( .IN1(n4240), .IN2(n5736), .QN(n4239) );
  OA22X1 U9239 ( .IN1(n5737), .IN2(n4253), .IN3(n4254), .IN4(n6047), .Q(g29291) );
  NAND2X0 U9240 ( .IN1(n4210), .IN2(n3289), .QN(n4253) );
  NOR2X0 U9241 ( .IN1(n4255), .IN2(n5737), .QN(n4254) );
  OA22X1 U9242 ( .IN1(n5738), .IN2(n4359), .IN3(n4360), .IN4(n6046), .Q(g29262) );
  NAND2X0 U9243 ( .IN1(n4210), .IN2(n3296), .QN(n4359) );
  NOR2X0 U9244 ( .IN1(n4361), .IN2(n5738), .QN(n4360) );
  OA22X1 U9245 ( .IN1(n5739), .IN2(n4207), .IN3(n4208), .IN4(n6046), .Q(g29309) );
  NAND2X0 U9246 ( .IN1(n4210), .IN2(n3295), .QN(n4207) );
  NOR2X0 U9247 ( .IN1(n4209), .IN2(n5739), .QN(n4208) );
  OA22X1 U9248 ( .IN1(n5740), .IN2(n4344), .IN3(n4345), .IN4(n6047), .Q(g29268) );
  NAND2X0 U9249 ( .IN1(n4210), .IN2(n3299), .QN(n4344) );
  NOR2X0 U9250 ( .IN1(n4346), .IN2(n5740), .QN(n4345) );
  OA22X1 U9251 ( .IN1(n5741), .IN2(n4223), .IN3(n4224), .IN4(n6047), .Q(g29303) );
  NAND2X0 U9252 ( .IN1(n4210), .IN2(n3292), .QN(n4223) );
  NOR2X0 U9253 ( .IN1(n4225), .IN2(n5741), .QN(n4224) );
  AO22X1 U9254 ( .IN1(g1373), .IN2(n3255), .IN3(n3256), .IN4(g1379), .Q(g33543) );
  NAND2X0 U9255 ( .IN1(n6218), .IN2(n3259), .QN(n3255) );
  OA21X1 U9256 ( .IN1(n3257), .IN2(n1572), .IN3(n6413), .Q(n3256) );
  OR3X1 U9257 ( .IN1(n3258), .IN2(g1379), .IN3(n1572), .Q(n3259) );
  AO22X1 U9258 ( .IN1(g1030), .IN2(n3263), .IN3(n3264), .IN4(g1036), .Q(g33541) );
  NAND2X0 U9259 ( .IN1(n6215), .IN2(n3267), .QN(n3263) );
  OA21X1 U9260 ( .IN1(n3265), .IN2(n1582), .IN3(n6411), .Q(n3264) );
  OR3X1 U9261 ( .IN1(n3266), .IN2(g1036), .IN3(n1582), .Q(n3267) );
  OA21X1 U9262 ( .IN1(n6117), .IN2(n1535), .IN3(g5694), .Q(g24343) );
  INVX0 U9263 ( .IN(n5153), .QN(n1535) );
  OA21X1 U9264 ( .IN1(n6116), .IN2(n1634), .IN3(g5348), .Q(g24339) );
  INVX0 U9265 ( .IN(n5158), .QN(n1634) );
  OA21X1 U9266 ( .IN1(n6117), .IN2(n1666), .IN3(g6386), .Q(g24351) );
  INVX0 U9267 ( .IN(n5143), .QN(n1666) );
  OA21X1 U9268 ( .IN1(n6116), .IN2(n1936), .IN3(g3343), .Q(g24270) );
  INVX0 U9269 ( .IN(n5190), .QN(n1936) );
  OA21X1 U9270 ( .IN1(n5117), .IN2(n5118), .IN3(n6369), .Q(g25609) );
  OA21X1 U9271 ( .IN1(n4818), .IN2(n5548), .IN3(test_so54), .Q(n5118) );
  OA21X1 U9272 ( .IN1(n4962), .IN2(n5287), .IN3(n2075), .Q(n5117) );
  OA21X1 U9273 ( .IN1(n6116), .IN2(n1523), .IN3(g6040), .Q(g24347) );
  INVX0 U9274 ( .IN(n5148), .QN(n1523) );
  OA21X1 U9275 ( .IN1(n6117), .IN2(n1675), .IN3(g6732), .Q(g24355) );
  INVX0 U9276 ( .IN(n5138), .QN(n1675) );
  OA21X1 U9277 ( .IN1(n6117), .IN2(n1503), .IN3(g4045), .Q(g24278) );
  INVX0 U9278 ( .IN(n5180), .QN(n1503) );
  OA21X1 U9279 ( .IN1(n6116), .IN2(n1707), .IN3(g3694), .Q(g24274) );
  INVX0 U9280 ( .IN(n5185), .QN(n1707) );
  OA21X1 U9281 ( .IN1(g5069), .IN2(n6118), .IN3(g5073), .Q(g25704) );
  OAI222X1 U9282 ( .IN1(n5309), .IN2(n2588), .IN3(n2586), .IN4(test_so99), 
        .IN5(n5391), .IN6(n6419), .QN(g34457) );
  NBUFFX2 U9283 ( .IN(g110), .Q(n6022) );
  NOR2X0 U9284 ( .IN1(g5073), .IN2(n6069), .QN(n5019) );
  NOR2X0 U9285 ( .IN1(n6083), .IN2(n5169), .QN(g24281) );
  XOR2X1 U9286 ( .IN1(g9251), .IN2(n5168), .Q(n5169) );
  NAND3X0 U9287 ( .IN1(n1469), .IN2(n5512), .IN3(g2208), .QN(n2998) );
  NAND3X0 U9288 ( .IN1(n3725), .IN2(n3463), .IN3(n3724), .QN(g31896) );
  NAND2X0 U9289 ( .IN1(g4477), .IN2(n6080), .QN(n3725) );
  NAND3X0 U9290 ( .IN1(n3457), .IN2(n3454), .IN3(n3461), .QN(g33041) );
  NAND2X0 U9291 ( .IN1(test_so56), .IN2(n6028), .QN(n3461) );
  NAND3X0 U9292 ( .IN1(n3723), .IN2(n3457), .IN3(n3724), .QN(g31897) );
  NAND2X0 U9293 ( .IN1(g4423), .IN2(n6080), .QN(n3723) );
  NAND3X0 U9294 ( .IN1(n3453), .IN2(n3454), .IN3(n3455), .QN(g33045) );
  NAND2X0 U9295 ( .IN1(g4567), .IN2(n6028), .QN(n3455) );
  NAND3X0 U9296 ( .IN1(n3462), .IN2(n3454), .IN3(n3465), .QN(g33038) );
  NAND2X0 U9297 ( .IN1(g4498), .IN2(n6028), .QN(n3465) );
  NAND3X0 U9298 ( .IN1(n3463), .IN2(n3454), .IN3(n3464), .QN(g33039) );
  NAND2X0 U9299 ( .IN1(g4501), .IN2(n6028), .QN(n3464) );
  NAND3X0 U9300 ( .IN1(n3463), .IN2(n3458), .IN3(n3466), .QN(g33037) );
  NAND2X0 U9301 ( .IN1(g4495), .IN2(n6027), .QN(n3466) );
  NAND3X0 U9302 ( .IN1(n3462), .IN2(n3458), .IN3(n3467), .QN(g33036) );
  NAND2X0 U9303 ( .IN1(g4480), .IN2(n6027), .QN(n3467) );
  NAND3X0 U9304 ( .IN1(n3453), .IN2(n3458), .IN3(n3460), .QN(g33042) );
  NAND2X0 U9305 ( .IN1(g4540), .IN2(n6028), .QN(n3460) );
  NAND3X0 U9306 ( .IN1(n3457), .IN2(n3458), .IN3(n3459), .QN(g33043) );
  NAND2X0 U9307 ( .IN1(test_so16), .IN2(n6028), .QN(n3459) );
  NOR3X0 U9308 ( .IN1(n2726), .IN2(g2599), .IN3(n5521), .QN(n2719) );
  NOR2X0 U9309 ( .IN1(n5022), .IN2(n5455), .QN(g25695) );
  OA221X1 U9310 ( .IN1(g5084), .IN2(g5073), .IN3(g5069), .IN4(n5681), .IN5(
        n6229), .Q(n5022) );
  AO222X1 U9311 ( .IN1(n5016), .IN2(n5753), .IN3(n5017), .IN4(g5097), .IN5(
        g5092), .IN6(n6108), .Q(g25698) );
  NOR2X0 U9312 ( .IN1(n5016), .IN2(n6063), .QN(n5017) );
  AO222X1 U9313 ( .IN1(n5014), .IN2(n5669), .IN3(n5015), .IN4(g20557), .IN5(
        g5097), .IN6(n6108), .Q(g25699) );
  NOR2X0 U9314 ( .IN1(n5014), .IN2(n6063), .QN(n5015) );
  ISOLANDX1 U9315 ( .D(n5016), .ISO(n5753), .Q(n5014) );
  NOR3X0 U9316 ( .IN1(n2727), .IN2(g2465), .IN3(n5522), .QN(n2720) );
  NOR2X0 U9317 ( .IN1(n5999), .IN2(n6000), .QN(n3174) );
  XOR2X1 U9318 ( .IN1(g490), .IN2(n6016), .Q(n5999) );
  XOR2X1 U9319 ( .IN1(g482), .IN2(n6018), .Q(n6000) );
  AO21X1 U9320 ( .IN1(g1996), .IN2(n2887), .IN3(n3193), .Q(g33568) );
  NOR4X0 U9321 ( .IN1(g2070), .IN2(n1292), .IN3(n3194), .IN4(n6117), .QN(n3193) );
  OA21X1 U9322 ( .IN1(g2040), .IN2(n1374), .IN3(n5355), .Q(n3194) );
  AO21X1 U9323 ( .IN1(g2153), .IN2(n2863), .IN3(n3172), .Q(g33576) );
  NOR4X0 U9324 ( .IN1(g2227), .IN2(n1293), .IN3(n3173), .IN4(n6118), .QN(n3172) );
  OA21X1 U9325 ( .IN1(g2197), .IN2(n2870), .IN3(n5356), .Q(n3173) );
  AO21X1 U9326 ( .IN1(test_so79), .IN2(n2817), .IN3(n3133), .Q(g33592) );
  NOR4X0 U9327 ( .IN1(g2495), .IN2(n3131), .IN3(n3134), .IN4(n6117), .QN(n3133) );
  OA21X1 U9328 ( .IN1(g2465), .IN2(n2824), .IN3(n5357), .Q(n3134) );
  NOR2X0 U9329 ( .IN1(n4878), .IN2(n6066), .QN(g26944) );
  NOR4X0 U9330 ( .IN1(n1390), .IN2(n4879), .IN3(n5298), .IN4(n4880), .QN(n4878) );
  NAND2X0 U9331 ( .IN1(g4358), .IN2(g4340), .QN(n4879) );
  NOR2X0 U9332 ( .IN1(n5212), .IN2(n6077), .QN(g24249) );
  OA22X1 U9333 ( .IN1(n5213), .IN2(n5850), .IN3(g1442), .IN4(n4475), .Q(n5212)
         );
  NOR2X0 U9334 ( .IN1(n4475), .IN2(n5617), .QN(n5213) );
  NOR2X0 U9335 ( .IN1(n5234), .IN2(n6077), .QN(g24233) );
  OA22X1 U9336 ( .IN1(n5235), .IN2(n5851), .IN3(test_so7), .IN4(n4499), .Q(
        n5234) );
  NOR2X0 U9337 ( .IN1(n4499), .IN2(n5618), .QN(n5235) );
  NOR2X0 U9338 ( .IN1(n2701), .IN2(n6077), .QN(g34253) );
  AND3X1 U9339 ( .IN1(g4462), .IN2(n2697), .IN3(test_so38), .Q(n2701) );
  NOR4X0 U9340 ( .IN1(n5189), .IN2(g16627), .IN3(g14451), .IN4(g16656), .QN(
        g24271) );
  AO221X1 U9341 ( .IN1(g16744), .IN2(n5699), .IN3(g13926), .IN4(n5433), .IN5(
        n6084), .Q(n5189) );
  NOR4X0 U9342 ( .IN1(n5142), .IN2(g17688), .IN3(g13099), .IN4(g17722), .QN(
        g24352) );
  AO221X1 U9343 ( .IN1(g17778), .IN2(n5700), .IN3(g14828), .IN4(n5434), .IN5(
        n6084), .Q(n5142) );
  NOR4X0 U9344 ( .IN1(n5184), .IN2(g16659), .IN3(g14518), .IN4(g16693), .QN(
        g24275) );
  AO221X1 U9345 ( .IN1(g16775), .IN2(n5701), .IN3(g13966), .IN4(n5435), .IN5(
        n6084), .Q(n5184) );
  NOR4X0 U9346 ( .IN1(n5194), .IN2(g16603), .IN3(g14421), .IN4(g16624), .QN(
        g24267) );
  AO221X1 U9347 ( .IN1(g16718), .IN2(n5702), .IN3(g13895), .IN4(n5436), .IN5(
        n6084), .Q(n5194) );
  NOR4X0 U9348 ( .IN1(n5147), .IN2(g17649), .IN3(g13085), .IN4(g17685), .QN(
        g24348) );
  AO221X1 U9349 ( .IN1(g17760), .IN2(n5703), .IN3(g14779), .IN4(n5437), .IN5(
        n6084), .Q(n5147) );
  NOR4X0 U9350 ( .IN1(n5162), .IN2(g17519), .IN3(g13039), .IN4(g17577), .QN(
        g24336) );
  AO221X1 U9351 ( .IN1(g17674), .IN2(n5704), .IN3(g14662), .IN4(n5438), .IN5(
        n6084), .Q(n5162) );
  NOR4X0 U9352 ( .IN1(n5157), .IN2(g17580), .IN3(g13049), .IN4(g17604), .QN(
        g24340) );
  AO221X1 U9353 ( .IN1(g17711), .IN2(n5705), .IN3(g14694), .IN4(n5439), .IN5(
        n6084), .Q(n5157) );
  OR2X1 U9354 ( .IN1(n5482), .IN2(g736), .Q(n4198) );
  NOR4X0 U9355 ( .IN1(g4871), .IN2(g4864), .IN3(g4836), .IN4(n1308), .QN(
        g34265) );
  NOR4X0 U9356 ( .IN1(g4681), .IN2(g4674), .IN3(g4646), .IN4(n1304), .QN(
        g34260) );
  NOR4X0 U9357 ( .IN1(n5229), .IN2(g17291), .IN3(g17400), .IN4(g17316), .QN(
        g24238) );
  AO21X1 U9358 ( .IN1(n5073), .IN2(n5230), .IN3(n6138), .Q(n5229) );
  NAND3X0 U9359 ( .IN1(n4194), .IN2(n5467), .IN3(n1986), .QN(n5230) );
  NOR4X0 U9360 ( .IN1(test_so68), .IN2(n4911), .IN3(n5059), .IN4(n6118), .QN(
        g25634) );
  AOI21X1 U9361 ( .IN1(n5060), .IN2(g12923), .IN3(g1395), .QN(n5059) );
  NOR4X0 U9362 ( .IN1(g979), .IN2(n4936), .IN3(n5083), .IN4(n6117), .QN(g25625) );
  AOI21X1 U9363 ( .IN1(n5084), .IN2(g12919), .IN3(g1052), .QN(n5083) );
  AO222X1 U9364 ( .IN1(n2887), .IN2(g2084), .IN3(n2888), .IN4(n2889), .IN5(
        g2070), .IN6(n6103), .Q(g33992) );
  NOR2X0 U9365 ( .IN1(n1374), .IN2(n6065), .QN(n2888) );
  XNOR2X1 U9366 ( .IN1(n2890), .IN2(n2891), .Q(n2889) );
  OA21X1 U9367 ( .IN1(g1996), .IN2(g2070), .IN3(g2084), .Q(n2890) );
  AO222X1 U9368 ( .IN1(n2817), .IN2(g2509), .IN3(n2818), .IN4(n2819), .IN5(
        g2495), .IN6(n6092), .Q(g34013) );
  NOR2X0 U9369 ( .IN1(n2824), .IN2(n6064), .QN(n2818) );
  XNOR2X1 U9370 ( .IN1(n2820), .IN2(n2821), .Q(n2819) );
  OA21X1 U9371 ( .IN1(test_so79), .IN2(g2495), .IN3(g2509), .Q(n2820) );
  AO222X1 U9372 ( .IN1(n2793), .IN2(g2643), .IN3(n2794), .IN4(n2795), .IN5(
        g2629), .IN6(n6093), .Q(g34020) );
  NOR2X0 U9373 ( .IN1(n2800), .IN2(n6064), .QN(n2794) );
  XNOR2X1 U9374 ( .IN1(n2796), .IN2(n2797), .Q(n2795) );
  OA21X1 U9375 ( .IN1(g2555), .IN2(g2629), .IN3(g2643), .Q(n2796) );
  AO222X1 U9376 ( .IN1(n2840), .IN2(g2375), .IN3(n2841), .IN4(n2842), .IN5(
        g2361), .IN6(n6091), .Q(g34006) );
  NOR2X0 U9377 ( .IN1(n2847), .IN2(n6064), .QN(n2841) );
  XNOR2X1 U9378 ( .IN1(n2843), .IN2(n2844), .Q(n2842) );
  OA21X1 U9379 ( .IN1(g2287), .IN2(g2361), .IN3(g2375), .Q(n2843) );
  AO222X1 U9380 ( .IN1(n2911), .IN2(g1950), .IN3(n2912), .IN4(n2913), .IN5(
        g1936), .IN6(n6101), .Q(g33985) );
  NOR2X0 U9381 ( .IN1(n1365), .IN2(n6065), .QN(n2912) );
  XNOR2X1 U9382 ( .IN1(n2914), .IN2(n2915), .Q(n2913) );
  OA21X1 U9383 ( .IN1(test_so8), .IN2(g1936), .IN3(g1950), .Q(n2914) );
  AO222X1 U9384 ( .IN1(n2863), .IN2(g2241), .IN3(n2864), .IN4(n2865), .IN5(
        g2227), .IN6(n6105), .Q(g33999) );
  NOR2X0 U9385 ( .IN1(n2870), .IN2(n6064), .QN(n2864) );
  XNOR2X1 U9386 ( .IN1(n2866), .IN2(n2867), .Q(n2865) );
  OA21X1 U9387 ( .IN1(g2153), .IN2(g2227), .IN3(g2241), .Q(n2866) );
  AO222X1 U9388 ( .IN1(n2957), .IN2(g1682), .IN3(n2958), .IN4(n2959), .IN5(
        g1668), .IN6(n6101), .Q(g33971) );
  NOR2X0 U9389 ( .IN1(n1347), .IN2(n6076), .QN(n2958) );
  XNOR2X1 U9390 ( .IN1(n2960), .IN2(n2961), .Q(n2959) );
  OA21X1 U9391 ( .IN1(g1592), .IN2(g1668), .IN3(g1682), .Q(n2960) );
  AND2X1 U9392 ( .IN1(n3726), .IN2(n3727), .Q(n3724) );
  NAND3X0 U9393 ( .IN1(n6415), .IN2(n5670), .IN3(g4372), .QN(n3727) );
  AO21X1 U9394 ( .IN1(n6016), .IN2(n6018), .IN3(n6028), .Q(n3726) );
  XNOR2X1 U9395 ( .IN1(g5084), .IN2(n5018), .Q(g25697) );
  NAND2X0 U9396 ( .IN1(g5092), .IN2(n6171), .QN(n5018) );
  XNOR2X1 U9397 ( .IN1(g990), .IN2(n5222), .Q(g24241) );
  NAND2X0 U9398 ( .IN1(n1740), .IN2(n6168), .QN(n5222) );
  XNOR2X1 U9399 ( .IN1(g1333), .IN2(n5200), .Q(g24257) );
  NAND2X0 U9400 ( .IN1(n1570), .IN2(n6154), .QN(n5200) );
  XNOR2X1 U9401 ( .IN1(g862), .IN2(n4942), .Q(g26910) );
  NAND2X0 U9402 ( .IN1(n6224), .IN2(n5305), .QN(n4942) );
  XNOR2X1 U9403 ( .IN1(g1430), .IN2(n5199), .Q(g24260) );
  NAND2X0 U9404 ( .IN1(g1548), .IN2(n6155), .QN(n5199) );
  XNOR2X1 U9405 ( .IN1(g1087), .IN2(n5221), .Q(g24244) );
  NAND2X0 U9406 ( .IN1(g1205), .IN2(n6166), .QN(n5221) );
  OAI221X1 U9407 ( .IN1(n3247), .IN2(n5758), .IN3(n3248), .IN4(n5412), .IN5(
        n3249), .QN(g33549) );
  NAND4X0 U9408 ( .IN1(n1349), .IN2(n6185), .IN3(n5417), .IN4(n5758), .QN(
        n3249) );
  OA21X1 U9409 ( .IN1(n3246), .IN2(n5417), .IN3(n6412), .Q(n3247) );
  OAI221X1 U9410 ( .IN1(n5030), .IN2(n5448), .IN3(n4331), .IN4(n5886), .IN5(
        n5031), .QN(g25683) );
  NAND4X0 U9411 ( .IN1(n1907), .IN2(n6182), .IN3(n5662), .IN4(n5448), .QN(
        n5031) );
  OA21X1 U9412 ( .IN1(n3298), .IN2(n5662), .IN3(n6363), .Q(n5030) );
  OAI221X1 U9413 ( .IN1(n4232), .IN2(n5747), .IN3(n4227), .IN4(n3761), .IN5(
        n4233), .QN(g29299) );
  NAND4X0 U9414 ( .IN1(g6159), .IN2(n4227), .IN3(n6173), .IN4(n5747), .QN(
        n4233) );
  OA21X1 U9415 ( .IN1(g6159), .IN2(n1566), .IN3(n6414), .Q(n4232) );
  OAI221X1 U9416 ( .IN1(n4997), .IN2(n5449), .IN3(n4240), .IN4(n5887), .IN5(
        n4998), .QN(g25735) );
  NAND4X0 U9417 ( .IN1(n1820), .IN2(n6183), .IN3(n5663), .IN4(n5449), .QN(
        n4998) );
  OA21X1 U9418 ( .IN1(n3294), .IN2(n5663), .IN3(n6362), .Q(n4997) );
  OAI221X1 U9419 ( .IN1(n3209), .IN2(n5450), .IN3(n3210), .IN4(n5845), .IN5(
        n3211), .QN(g33565) );
  NAND4X0 U9420 ( .IN1(n1367), .IN2(n6188), .IN3(n5664), .IN4(n5450), .QN(
        n3211) );
  OA21X1 U9421 ( .IN1(n3208), .IN2(n5664), .IN3(n6371), .Q(n3209) );
  OAI221X1 U9422 ( .IN1(n3108), .IN2(n5759), .IN3(n3109), .IN4(n5278), .IN5(
        n3110), .QN(g33605) );
  NAND4X0 U9423 ( .IN1(n1335), .IN2(n6180), .IN3(n5418), .IN4(n5759), .QN(
        n3110) );
  OA21X1 U9424 ( .IN1(n3107), .IN2(n5418), .IN3(n6368), .Q(n3108) );
  OAI221X1 U9425 ( .IN1(n4217), .IN2(n5748), .IN3(n4212), .IN4(n2474), .IN5(
        n4218), .QN(g29305) );
  NAND4X0 U9426 ( .IN1(g6505), .IN2(n4212), .IN3(n6168), .IN4(n5748), .QN(
        n4218) );
  OA21X1 U9427 ( .IN1(g6505), .IN2(n1674), .IN3(n6410), .Q(n4217) );
  OAI221X1 U9428 ( .IN1(n3168), .IN2(n5760), .IN3(n3169), .IN4(n5410), .IN5(
        n3170), .QN(g33581) );
  NAND4X0 U9429 ( .IN1(n1311), .IN2(n6189), .IN3(n5419), .IN4(n5760), .QN(
        n3170) );
  OA21X1 U9430 ( .IN1(n3167), .IN2(n5419), .IN3(n6371), .Q(n3168) );
  OAI221X1 U9431 ( .IN1(n3229), .IN2(n5451), .IN3(n3230), .IN4(n5847), .IN5(
        n3231), .QN(g33557) );
  NAND4X0 U9432 ( .IN1(n1358), .IN2(n6187), .IN3(n5665), .IN4(n5451), .QN(
        n3231) );
  OA21X1 U9433 ( .IN1(n3228), .IN2(n5665), .IN3(n6412), .Q(n3229) );
  OAI221X1 U9434 ( .IN1(n4247), .IN2(n5749), .IN3(n4242), .IN4(n3760), .IN5(
        n4248), .QN(g29293) );
  NAND4X0 U9435 ( .IN1(g5813), .IN2(n4242), .IN3(n6172), .IN4(n5749), .QN(
        n4248) );
  OA21X1 U9436 ( .IN1(g5813), .IN2(n1563), .IN3(n6412), .Q(n4247) );
  OAI221X1 U9437 ( .IN1(n3128), .IN2(n5761), .IN3(n3129), .IN4(n5411), .IN5(
        n3130), .QN(g33597) );
  NAND4X0 U9438 ( .IN1(n1327), .IN2(n6184), .IN3(n5420), .IN4(n5761), .QN(
        n3130) );
  OA21X1 U9439 ( .IN1(n3127), .IN2(n5420), .IN3(n6367), .Q(n3128) );
  OAI221X1 U9440 ( .IN1(n3149), .IN2(n5762), .IN3(n3150), .IN4(n5279), .IN5(
        n3151), .QN(g33589) );
  NAND4X0 U9441 ( .IN1(n1319), .IN2(n6194), .IN3(n5421), .IN4(n5762), .QN(
        n3151) );
  OA21X1 U9442 ( .IN1(n3148), .IN2(n5421), .IN3(n6370), .Q(n3149) );
  OAI221X1 U9443 ( .IN1(n3189), .IN2(n5452), .IN3(n3190), .IN4(n5848), .IN5(
        n3191), .QN(g33573) );
  NAND4X0 U9444 ( .IN1(n1376), .IN2(n6193), .IN3(n5666), .IN4(n5452), .QN(
        n3191) );
  OA21X1 U9445 ( .IN1(n3188), .IN2(n5666), .IN3(n6370), .Q(n3189) );
  OAI221X1 U9446 ( .IN1(n4992), .IN2(n5453), .IN3(n4225), .IN4(n5888), .IN5(
        n4993), .QN(g25749) );
  NAND4X0 U9447 ( .IN1(n1513), .IN2(n6192), .IN3(n5667), .IN4(n5453), .QN(
        n4993) );
  OA21X1 U9448 ( .IN1(n3292), .IN2(n5667), .IN3(n6359), .Q(n4992) );
  OAI221X1 U9449 ( .IN1(n5035), .IN2(n5454), .IN3(n4346), .IN4(n5889), .IN5(
        n5036), .QN(g25669) );
  NAND4X0 U9450 ( .IN1(n1679), .IN2(n6181), .IN3(n5668), .IN4(n5454), .QN(
        n5036) );
  OA21X1 U9451 ( .IN1(n3299), .IN2(n5668), .IN3(n6362), .Q(n5035) );
  OAI221X1 U9452 ( .IN1(n3063), .IN2(g4104), .IN3(n5715), .IN4(n6267), .IN5(
        n3064), .QN(g33615) );
  ISOLANDX1 U9453 ( .D(n3065), .ISO(n1437), .Q(n3064) );
  NAND3X0 U9454 ( .IN1(n6415), .IN2(n3063), .IN3(g4104), .QN(n3065) );
  NAND2X0 U9455 ( .IN1(n1645), .IN2(g4108), .QN(n3063) );
  NAND2X0 U9456 ( .IN1(g4575), .IN2(n1402), .QN(n3457) );
  XOR2X1 U9457 ( .IN1(DFF_228_n1), .IN2(n4857), .Q(g26965) );
  NAND2X0 U9458 ( .IN1(g10306), .IN2(n6161), .QN(n4857) );
  NOR3X0 U9459 ( .IN1(g358), .IN2(g8719), .IN3(n6082), .QN(g25595) );
  NOR3X0 U9460 ( .IN1(n4203), .IN2(n5250), .IN3(n6081), .QN(g24210) );
  OA22X1 U9461 ( .IN1(n5251), .IN2(n5306), .IN3(n5402), .IN4(n5606), .Q(n5250)
         );
  NOR2X0 U9462 ( .IN1(g168), .IN2(g174), .QN(n5251) );
  NAND4X0 U9463 ( .IN1(n6195), .IN2(n2699), .IN3(n2697), .IN4(n5671), .QN(
        g34255) );
  NAND2X0 U9464 ( .IN1(test_so38), .IN2(g4473), .QN(n2699) );
  AO22X1 U9465 ( .IN1(n6136), .IN2(g1740), .IN3(n2951), .IN4(n6284), .Q(g33973) );
  OAI22X1 U9466 ( .IN1(n2933), .IN2(n2952), .IN3(n1359), .IN4(n5817), .QN(
        n2951) );
  INVX0 U9467 ( .IN(n2952), .QN(n1359) );
  NAND3X0 U9468 ( .IN1(n2953), .IN2(n5504), .IN3(g1728), .QN(n2952) );
  AOI21X1 U9469 ( .IN1(n4055), .IN2(n4056), .IN3(n6122), .QN(n4044) );
  NAND4X0 U9470 ( .IN1(n4059), .IN2(n4060), .IN3(n4061), .IN4(n4050), .QN(
        n4055) );
  AO221X1 U9471 ( .IN1(n2140), .IN2(g2783), .IN3(n2138), .IN4(g2787), .IN5(
        n4057), .Q(n4056) );
  OR2X1 U9472 ( .IN1(n4052), .IN2(g2079), .Q(n4060) );
  AOI21X1 U9473 ( .IN1(n4045), .IN2(n4046), .IN3(n6122), .QN(n4043) );
  NAND4X0 U9474 ( .IN1(n4047), .IN2(n4048), .IN3(n4049), .IN4(n4050), .QN(
        n4046) );
  AO221X1 U9475 ( .IN1(n2140), .IN2(g2815), .IN3(n2138), .IN4(g2819), .IN5(
        n4053), .Q(n4045) );
  OR2X1 U9476 ( .IN1(n4052), .IN2(g2638), .Q(n4048) );
  OAI22X1 U9477 ( .IN1(n1297), .IN2(n5391), .IN3(n2578), .IN4(n5727), .QN(
        g34460) );
  OA21X1 U9478 ( .IN1(test_so3), .IN2(n2579), .IN3(n6364), .Q(n2578) );
  OAI22X1 U9479 ( .IN1(n6322), .IN2(n5348), .IN3(n5165), .IN4(n5166), .QN(
        g24334) );
  NAND4X0 U9480 ( .IN1(n5303), .IN2(n5365), .IN3(n5274), .IN4(n5608), .QN(
        n5165) );
  NAND4X0 U9481 ( .IN1(n5164), .IN2(n1532), .IN3(g4340), .IN4(n5539), .QN(
        n5166) );
  OAI22X1 U9482 ( .IN1(n2564), .IN2(n5283), .IN3(n1308), .IN4(n2565), .QN(
        g34466) );
  NAND2X0 U9483 ( .IN1(g4843), .IN2(n5283), .QN(n2565) );
  OA21X1 U9484 ( .IN1(g4843), .IN2(n2560), .IN3(n6366), .Q(n2564) );
  OAI22X1 U9485 ( .IN1(n6138), .IN2(g218), .IN3(n5595), .IN4(n6352), .QN(
        g25591) );
  OAI22X1 U9486 ( .IN1(n2574), .IN2(n5656), .IN3(n1304), .IN4(n2575), .QN(
        g34462) );
  NAND2X0 U9487 ( .IN1(test_so19), .IN2(n5656), .QN(n2575) );
  OA21X1 U9488 ( .IN1(test_so19), .IN2(n2570), .IN3(n6365), .Q(n2574) );
  OAI22X1 U9489 ( .IN1(n6304), .IN2(n5653), .IN3(n1299), .IN4(n2694), .QN(
        g34257) );
  OA22X1 U9490 ( .IN1(n5298), .IN2(n2695), .IN3(test_so81), .IN4(n2693), .Q(
        n2694) );
  NAND2X0 U9491 ( .IN1(n6188), .IN2(n2693), .QN(n2695) );
  OAI22X1 U9492 ( .IN1(n6304), .IN2(n5298), .IN3(n1299), .IN4(n2691), .QN(
        g34258) );
  OA22X1 U9493 ( .IN1(n5348), .IN2(n2692), .IN3(g4358), .IN4(n2609), .Q(n2691)
         );
  NAND2X0 U9494 ( .IN1(n6665), .IN2(n2609), .QN(n2692) );
  OAI22X1 U9495 ( .IN1(n4125), .IN2(n6146), .IN3(n4126), .IN4(n5783), .QN(
        g30362) );
  OA22X1 U9496 ( .IN1(n4127), .IN2(n4128), .IN3(n1612), .IN4(n5890), .Q(n4125)
         );
  OA21X1 U9497 ( .IN1(n5462), .IN2(n4127), .IN3(n6407), .Q(n4126) );
  OAI22X1 U9498 ( .IN1(n5383), .IN2(n3486), .IN3(n3487), .IN4(n5645), .QN(
        g33028) );
  OA21X1 U9499 ( .IN1(g3522), .IN2(n1281), .IN3(n6409), .Q(n3487) );
  OAI22X1 U9500 ( .IN1(n5386), .IN2(n3401), .IN3(n3402), .IN4(n5646), .QN(
        g33069) );
  OA21X1 U9501 ( .IN1(g6565), .IN2(n1283), .IN3(n6413), .Q(n3402) );
  OAI22X1 U9502 ( .IN1(n5389), .IN2(n3431), .IN3(n3432), .IN4(n5647), .QN(
        g33054) );
  OA21X1 U9503 ( .IN1(g5527), .IN2(n1285), .IN3(n6411), .Q(n3432) );
  OAI22X1 U9504 ( .IN1(n5387), .IN2(n3476), .IN3(n3477), .IN4(n5648), .QN(
        g33033) );
  OA21X1 U9505 ( .IN1(g3873), .IN2(n1282), .IN3(n6408), .Q(n3477) );
  OAI22X1 U9506 ( .IN1(n5388), .IN2(n3421), .IN3(n3422), .IN4(n5649), .QN(
        g33059) );
  OA21X1 U9507 ( .IN1(g5873), .IN2(n1286), .IN3(n6411), .Q(n3422) );
  OAI22X1 U9508 ( .IN1(n5384), .IN2(n3441), .IN3(n3442), .IN4(n5650), .QN(
        g33049) );
  OA21X1 U9509 ( .IN1(g5180), .IN2(n1284), .IN3(n6410), .Q(n3442) );
  OAI22X1 U9510 ( .IN1(n5385), .IN2(n3411), .IN3(n3412), .IN4(n5651), .QN(
        g33064) );
  OA21X1 U9511 ( .IN1(g6219), .IN2(n1287), .IN3(n6406), .Q(n3412) );
  OAI22X1 U9512 ( .IN1(n6319), .IN2(n5328), .IN3(n4491), .IN4(n6141), .QN(
        g29234) );
  OA22X1 U9513 ( .IN1(n4492), .IN2(n4493), .IN3(n4494), .IN4(n5864), .Q(n4491)
         );
  NAND2X0 U9514 ( .IN1(n4496), .IN2(n4495), .QN(n4493) );
  OAI22X1 U9515 ( .IN1(n5028), .IN2(n5416), .IN3(n5027), .IN4(n5029), .QN(
        g25686) );
  NAND2X0 U9516 ( .IN1(g4057), .IN2(n5416), .QN(n5029) );
  OA21X1 U9517 ( .IN1(g4057), .IN2(n5729), .IN3(n6361), .Q(n5028) );
  OAI22X1 U9518 ( .IN1(n6138), .IN2(g4239), .IN3(n5764), .IN4(n6353), .QN(
        g21892) );
  OAI22X1 U9519 ( .IN1(n4113), .IN2(n6145), .IN3(n4114), .IN4(n5784), .QN(
        g30367) );
  OA22X1 U9520 ( .IN1(n4115), .IN2(n4116), .IN3(n1856), .IN4(n5891), .Q(n4113)
         );
  OA21X1 U9521 ( .IN1(n5463), .IN2(n4115), .IN3(n6407), .Q(n4114) );
  OAI22X1 U9522 ( .IN1(n4137), .IN2(n6145), .IN3(n4138), .IN4(n5785), .QN(
        g30357) );
  OA21X1 U9523 ( .IN1(n5464), .IN2(n4139), .IN3(n6409), .Q(n4138) );
  OA22X1 U9524 ( .IN1(n4139), .IN2(n4140), .IN3(n1852), .IN4(n5892), .Q(n4137)
         );
  OAI22X1 U9525 ( .IN1(n4349), .IN2(n6145), .IN3(n4350), .IN4(n5786), .QN(
        g29266) );
  OA22X1 U9526 ( .IN1(n1594), .IN2(n4351), .IN3(n4348), .IN4(n5868), .Q(n4349)
         );
  OA21X1 U9527 ( .IN1(n1594), .IN2(n5424), .IN3(n6365), .Q(n4350) );
  OAI22X1 U9528 ( .IN1(n6319), .IN2(n5290), .IN3(n4474), .IN4(n6141), .QN(
        g29238) );
  OA22X1 U9529 ( .IN1(n4475), .IN2(n4476), .IN3(n4477), .IN4(n5865), .Q(n4474)
         );
  NAND2X0 U9530 ( .IN1(n4472), .IN2(n4478), .QN(n4476) );
  OAI22X1 U9531 ( .IN1(n6320), .IN2(n5289), .IN3(n4467), .IN4(n6140), .QN(
        g29239) );
  OA22X1 U9532 ( .IN1(n4468), .IN2(n4469), .IN3(n4470), .IN4(n5866), .Q(n4467)
         );
  NAND2X0 U9533 ( .IN1(n4472), .IN2(n4471), .QN(n4469) );
  OAI22X1 U9534 ( .IN1(n6323), .IN2(n5657), .IN3(n4817), .IN4(n6142), .QN(
        g28048) );
  OA22X1 U9535 ( .IN1(n4818), .IN2(n4819), .IN3(n4820), .IN4(n5520), .Q(n4817)
         );
  OA21X1 U9536 ( .IN1(test_so70), .IN2(n5821), .IN3(n2075), .Q(n4820) );
  OAI22X1 U9537 ( .IN1(n6321), .IN2(n5733), .IN3(n4520), .IN4(n5101), .QN(
        g25617) );
  OA22X1 U9538 ( .IN1(g817), .IN2(n5102), .IN3(n5822), .IN4(n4545), .Q(n5101)
         );
  OAI22X1 U9539 ( .IN1(n6323), .IN2(n5305), .IN3(n4943), .IN4(n6140), .QN(
        g26909) );
  OA22X1 U9540 ( .IN1(g896), .IN2(n5682), .IN3(g890), .IN4(n5431), .Q(n4943)
         );
  OAI22X1 U9541 ( .IN1(n4258), .IN2(n5805), .IN3(n4259), .IN4(n6140), .QN(
        g29289) );
  OA22X1 U9542 ( .IN1(n1561), .IN2(n4260), .IN3(n4257), .IN4(n5869), .Q(n4259)
         );
  OA21X1 U9543 ( .IN1(n1561), .IN2(n5425), .IN3(n6371), .Q(n4258) );
  OAI22X1 U9544 ( .IN1(n3746), .IN2(n5695), .IN3(n2709), .IN4(n3747), .QN(
        g31865) );
  NAND2X0 U9545 ( .IN1(test_so51), .IN2(n5695), .QN(n3747) );
  OA21X1 U9546 ( .IN1(test_so51), .IN2(n3748), .IN3(n6404), .Q(n3746) );
  OAI22X1 U9547 ( .IN1(n4213), .IN2(n5806), .IN3(n4214), .IN4(n6140), .QN(
        g29307) );
  OA22X1 U9548 ( .IN1(n1674), .IN2(n4215), .IN3(n4212), .IN4(n5870), .Q(n4214)
         );
  OA21X1 U9549 ( .IN1(n1674), .IN2(n5426), .IN3(n6413), .Q(n4213) );
  OAI22X1 U9550 ( .IN1(n4273), .IN2(n5807), .IN3(n4274), .IN4(n6140), .QN(
        g29283) );
  OA22X1 U9551 ( .IN1(n1559), .IN2(n4275), .IN3(n4272), .IN4(n5871), .Q(n4274)
         );
  OA21X1 U9552 ( .IN1(n1559), .IN2(n5427), .IN3(n6369), .Q(n4273) );
  OAI22X1 U9553 ( .IN1(n4334), .IN2(n5808), .IN3(n4335), .IN4(n6140), .QN(
        g29272) );
  OA22X1 U9554 ( .IN1(n1502), .IN2(n4336), .IN3(n4333), .IN4(n5872), .Q(n4335)
         );
  OA21X1 U9555 ( .IN1(n1502), .IN2(n5428), .IN3(n6369), .Q(n4334) );
  OAI22X1 U9556 ( .IN1(n4243), .IN2(n5809), .IN3(n4244), .IN4(n6140), .QN(
        g29295) );
  OA22X1 U9557 ( .IN1(n1563), .IN2(n4245), .IN3(n4242), .IN4(n5873), .Q(n4244)
         );
  OA21X1 U9558 ( .IN1(n1563), .IN2(n5429), .IN3(n6414), .Q(n4243) );
  OAI22X1 U9559 ( .IN1(n4228), .IN2(n5810), .IN3(n4229), .IN4(n6140), .QN(
        g29301) );
  OA22X1 U9560 ( .IN1(n1566), .IN2(n4230), .IN3(n4227), .IN4(n5874), .Q(n4229)
         );
  OA21X1 U9561 ( .IN1(n1566), .IN2(n5430), .IN3(n6408), .Q(n4228) );
  OAI22X1 U9562 ( .IN1(n6321), .IN2(n5796), .IN3(n5209), .IN4(n6140), .QN(
        g24253) );
  AOI22X1 U9563 ( .IN1(n5302), .IN2(g1532), .IN3(g1521), .IN4(n6024), .QN(
        n5209) );
  OAI22X1 U9564 ( .IN1(n6304), .IN2(n5771), .IN3(n2685), .IN4(n6141), .QN(
        g34261) );
  OA22X1 U9565 ( .IN1(n5862), .IN2(n2686), .IN3(n2687), .IN4(n1380), .Q(n2685)
         );
  INVX0 U9566 ( .IN(n2686), .QN(n1380) );
  OAI22X1 U9567 ( .IN1(n6301), .IN2(n5772), .IN3(n2656), .IN4(n6141), .QN(
        g34268) );
  OA22X1 U9568 ( .IN1(n5875), .IN2(n2657), .IN3(n2658), .IN4(n1388), .Q(n2656)
         );
  INVX0 U9569 ( .IN(n2657), .QN(n1388) );
  OAI22X1 U9570 ( .IN1(n6302), .IN2(n5773), .IN3(n2681), .IN4(n6142), .QN(
        g34262) );
  OA22X1 U9571 ( .IN1(n5876), .IN2(n2682), .IN3(n2683), .IN4(n1382), .Q(n2681)
         );
  INVX0 U9572 ( .IN(n2682), .QN(n1382) );
  OAI22X1 U9573 ( .IN1(n6301), .IN2(n5774), .IN3(n2664), .IN4(n6142), .QN(
        g34266) );
  OA22X1 U9574 ( .IN1(n5863), .IN2(n2665), .IN3(n2666), .IN4(n1385), .Q(n2664)
         );
  INVX0 U9575 ( .IN(n2665), .QN(n1385) );
  OAI22X1 U9576 ( .IN1(n6302), .IN2(n5775), .IN3(n2677), .IN4(n6141), .QN(
        g34263) );
  OA22X1 U9577 ( .IN1(n5877), .IN2(n2678), .IN3(n2679), .IN4(n1383), .Q(n2677)
         );
  INVX0 U9578 ( .IN(n2678), .QN(n1383) );
  OAI22X1 U9579 ( .IN1(n6303), .IN2(n5776), .IN3(n2660), .IN4(n6141), .QN(
        g34267) );
  OA22X1 U9580 ( .IN1(n5878), .IN2(n2661), .IN3(n2662), .IN4(n1387), .Q(n2660)
         );
  INVX0 U9581 ( .IN(n2661), .QN(n1387) );
  OAI22X1 U9582 ( .IN1(n6319), .IN2(n5630), .IN3(n5231), .IN4(n6140), .QN(
        g24237) );
  AOI22X1 U9583 ( .IN1(n5304), .IN2(g1189), .IN3(g1178), .IN4(n6021), .QN(
        n5231) );
  OAI22X1 U9584 ( .IN1(n5080), .IN2(n5691), .IN3(n5081), .IN4(n5341), .QN(
        g25626) );
  OA221X1 U9585 ( .IN1(n1695), .IN2(n5341), .IN3(n4924), .IN4(n5082), .IN5(
        n6571), .Q(n5080) );
  OA22X1 U9586 ( .IN1(n1606), .IN2(n5691), .IN3(g1141), .IN4(n6137), .Q(n5081)
         );
  NAND2X0 U9587 ( .IN1(n1695), .IN2(n5341), .QN(n5082) );
  OAI22X1 U9588 ( .IN1(n4926), .IN2(n5692), .IN3(n4927), .IN4(n5329), .QN(
        g26916) );
  OA221X1 U9589 ( .IN1(n1693), .IN2(n5329), .IN3(n4924), .IN4(n4928), .IN5(
        n6232), .Q(n4926) );
  OA22X1 U9590 ( .IN1(n1606), .IN2(n5692), .IN3(g1124), .IN4(n6137), .Q(n4927)
         );
  NAND2X0 U9591 ( .IN1(n1693), .IN2(n5329), .QN(n4928) );
  OAI22X1 U9592 ( .IN1(n4897), .IN2(n5696), .IN3(n4898), .IN4(n5289), .QN(
        g26924) );
  OA221X1 U9593 ( .IN1(n1775), .IN2(n5289), .IN3(n4899), .IN4(n4900), .IN5(
        n6231), .Q(n4897) );
  OA22X1 U9594 ( .IN1(n1655), .IN2(n5696), .IN3(g1437), .IN4(n6137), .Q(n4898)
         );
  NAND2X0 U9595 ( .IN1(n1775), .IN2(n5289), .QN(n4900) );
  OAI22X1 U9596 ( .IN1(n4901), .IN2(n5693), .IN3(n4902), .IN4(n5290), .QN(
        g26923) );
  OA221X1 U9597 ( .IN1(n1776), .IN2(n5290), .IN3(n4899), .IN4(n4903), .IN5(
        n6665), .Q(n4901) );
  OA22X1 U9598 ( .IN1(n1655), .IN2(n5693), .IN3(g1467), .IN4(n6137), .Q(n4902)
         );
  NAND2X0 U9599 ( .IN1(n1776), .IN2(n5290), .QN(n4903) );
  OAI22X1 U9600 ( .IN1(n4922), .IN2(n5697), .IN3(n4923), .IN4(n5328), .QN(
        g26917) );
  OA221X1 U9601 ( .IN1(n1692), .IN2(n5328), .IN3(n4924), .IN4(n4925), .IN5(
        n6665), .Q(n4922) );
  OA22X1 U9602 ( .IN1(n1606), .IN2(n5697), .IN3(g1094), .IN4(n6137), .Q(n4923)
         );
  NAND2X0 U9603 ( .IN1(n1692), .IN2(n5328), .QN(n4925) );
  OAI22X1 U9604 ( .IN1(n6320), .IN2(n5766), .IN3(n4975), .IN4(n6143), .QN(
        g26884) );
  OA21X1 U9605 ( .IN1(n4971), .IN2(n4976), .IN3(n4977), .Q(n4975) );
  NAND4X0 U9606 ( .IN1(n5282), .IN2(n5317), .IN3(n5456), .IN4(n5766), .QN(
        n4977) );
  OA221X1 U9607 ( .IN1(g336), .IN2(n5317), .IN3(n5282), .IN4(n5824), .IN5(
        n5456), .Q(n4976) );
  OAI22X1 U9608 ( .IN1(n6318), .IN2(n5587), .IN3(n2970), .IN4(n6144), .QN(
        g33968) );
  OA22X1 U9609 ( .IN1(n2956), .IN2(n2971), .IN3(n1344), .IN4(n5855), .Q(n2970)
         );
  INVX0 U9610 ( .IN(n2971), .QN(n1344) );
  OAI22X1 U9611 ( .IN1(n6308), .IN2(n5685), .IN3(n2831), .IN4(n6142), .QN(
        g34010) );
  OA22X1 U9612 ( .IN1(n2816), .IN2(n2832), .IN3(n1332), .IN4(n5856), .Q(n2831)
         );
  INVX0 U9613 ( .IN(n2832), .QN(n1332) );
  NAND2X0 U9614 ( .IN1(n4969), .IN2(n4970), .QN(g26889) );
  NAND4X0 U9615 ( .IN1(g329), .IN2(n4971), .IN3(n6170), .IN4(DFF_709_n1), .QN(
        n4970) );
  NAND2X0 U9616 ( .IN1(g20763), .IN2(n6080), .QN(n4969) );
  OA221X1 U9617 ( .IN1(n3311), .IN2(n5492), .IN3(n3312), .IN4(n5333), .IN5(
        n3336), .Q(n3335) );
  AOI222X1 U9618 ( .IN1(n1791), .IN2(g554), .IN3(n1795), .IN4(g582), .IN5(
        n1794), .IN6(g622), .QN(n3336) );
  AOI222X1 U9619 ( .IN1(n1793), .IN2(g2878), .IN3(n2459), .IN4(g2965), .IN5(
        n6001), .IN6(test_so22), .QN(n3371) );
  AOI221X1 U9620 ( .IN1(n1793), .IN2(g2848), .IN3(n6001), .IN4(test_so1), 
        .IN5(n3316), .QN(n3308) );
  AO22X1 U9621 ( .IN1(n2546), .IN2(g2844), .IN3(n2459), .IN4(g2902), .Q(n3316)
         );
  NAND2X0 U9622 ( .IN1(n4711), .IN2(n4712), .QN(g28082) );
  NAND3X0 U9623 ( .IN1(n6414), .IN2(n5752), .IN3(n2417), .QN(n4712) );
  OAI21X1 U9624 ( .IN1(n4713), .IN2(n6139), .IN3(g4521), .QN(n4711) );
  NAND2X0 U9625 ( .IN1(n2780), .IN2(n2781), .QN(g34023) );
  AO21X1 U9626 ( .IN1(n6202), .IN2(n2783), .IN3(DFF_491_n1), .Q(n2780) );
  NAND3X0 U9627 ( .IN1(n2778), .IN2(n2782), .IN3(n6325), .QN(n2781) );
  NAND4X0 U9628 ( .IN1(g4561), .IN2(g4558), .IN3(g4555), .IN4(n2782), .QN(
        n2783) );
  AOI21X1 U9629 ( .IN1(g847), .IN2(g843), .IN3(n6122), .QN(n4951) );
  AND3X1 U9630 ( .IN1(n3381), .IN2(g28), .IN3(n3382), .Q(n6001) );
  OAI22X1 U9631 ( .IN1(n6311), .IN2(n5688), .IN3(n2877), .IN4(n6142), .QN(
        g33996) );
  OA22X1 U9632 ( .IN1(n2862), .IN2(n2878), .IN3(n1316), .IN4(n5857), .Q(n2877)
         );
  INVX0 U9633 ( .IN(n2878), .QN(n1316) );
  OAI22X1 U9634 ( .IN1(n6307), .IN2(n5684), .IN3(n2807), .IN4(n6141), .QN(
        g34017) );
  OA22X1 U9635 ( .IN1(n2792), .IN2(n2808), .IN3(n1340), .IN4(n5858), .Q(n2807)
         );
  INVX0 U9636 ( .IN(n2808), .QN(n1340) );
  OAI22X1 U9637 ( .IN1(n6310), .IN2(n5687), .IN3(n2854), .IN4(n6142), .QN(
        g34003) );
  OA22X1 U9638 ( .IN1(n2839), .IN2(n2855), .IN3(n1324), .IN4(n5859), .Q(n2854)
         );
  INVX0 U9639 ( .IN(n2855), .QN(n1324) );
  AO22X1 U9640 ( .IN1(n6134), .IN2(g2008), .IN3(n2904), .IN4(n6289), .Q(g33987) );
  OAI22X1 U9641 ( .IN1(n2886), .IN2(n2905), .IN3(n1377), .IN4(n5818), .QN(
        n2904) );
  INVX0 U9642 ( .IN(n2905), .QN(n1377) );
  NAND3X0 U9643 ( .IN1(n2906), .IN2(n5505), .IN3(g1996), .QN(n2905) );
  OA21X1 U9644 ( .IN1(n4321), .IN2(n4698), .IN3(g4646), .Q(g28753) );
  OA21X1 U9645 ( .IN1(n5363), .IN2(n3196), .IN3(g17291), .Q(g27831) );
  NAND4X0 U9646 ( .IN1(g8403), .IN2(g8283), .IN3(n2668), .IN4(n1591), .QN(
        g33935) );
  INVX0 U9647 ( .IN(g34649), .QN(n1591) );
  NAND4X0 U9648 ( .IN1(g8353), .IN2(g8235), .IN3(n2668), .IN4(n1686), .QN(
        g33636) );
  INVX0 U9649 ( .IN(g34657), .QN(n1686) );
  NAND4X0 U9650 ( .IN1(n4298), .IN2(n4299), .IN3(n4300), .IN4(n4301), .QN(
        g34649) );
  NAND2X0 U9651 ( .IN1(g4955), .IN2(n2134), .QN(n4298) );
  NAND4X0 U9652 ( .IN1(n4320), .IN2(n4321), .IN3(n4322), .IN4(n4323), .QN(
        g34657) );
  NAND2X0 U9653 ( .IN1(g4765), .IN2(n2102), .QN(n4320) );
  AOI21X1 U9654 ( .IN1(n3195), .IN2(g479), .IN3(n5305), .QN(g33894) );
  NOR4X0 U9655 ( .IN1(n5481), .IN2(n4828), .IN3(n2076), .IN4(g504), .QN(n4532)
         );
  NAND2X0 U9656 ( .IN1(g24174), .IN2(g2873), .QN(g34436) );
  NAND2X0 U9657 ( .IN1(g24174), .IN2(g2868), .QN(g34437) );
  NAND4X0 U9658 ( .IN1(n1986), .IN2(n5227), .IN3(n4194), .IN4(n5467), .QN(
        n5226) );
  XNOR2X1 U9659 ( .IN1(n5320), .IN2(g1236), .Q(n5227) );
  NAND4X0 U9660 ( .IN1(n1571), .IN2(n5205), .IN3(n4176), .IN4(n5466), .QN(
        n5204) );
  XNOR2X1 U9661 ( .IN1(g1579), .IN2(n5319), .Q(n5205) );
  AO21X1 U9662 ( .IN1(n1490), .IN2(n1300), .IN3(DFF_961_n1), .Q(n2582) );
  OA221X1 U9663 ( .IN1(n2632), .IN2(n5609), .IN3(n5404), .IN4(n2637), .IN5(
        n5137), .Q(g33079) );
  AO221X1 U9664 ( .IN1(n5301), .IN2(n5545), .IN3(g2724), .IN4(n5379), .IN5(
        g2729), .Q(n5137) );
  OA221X1 U9665 ( .IN1(n2632), .IN2(n5610), .IN3(n2637), .IN4(n5403), .IN5(
        n5136), .Q(g33435) );
  AO221X1 U9666 ( .IN1(n5301), .IN2(n5544), .IN3(g2724), .IN4(n5378), .IN5(
        g2729), .Q(n5136) );
  NAND2X0 U9667 ( .IN1(g3179), .IN2(n5603), .QN(n3495) );
  NAND2X0 U9668 ( .IN1(g13259), .IN2(n1694), .QN(n4504) );
  NAND2X0 U9669 ( .IN1(g13272), .IN2(n2035), .QN(n4480) );
  NAND2X0 U9670 ( .IN1(g4688), .IN2(n4697), .QN(n3027) );
  OR3X1 U9671 ( .IN1(n5613), .IN2(n4326), .IN3(n4698), .Q(n4697) );
  NAND2X0 U9672 ( .IN1(g4878), .IN2(n4752), .QN(n3069) );
  OR3X1 U9673 ( .IN1(n5614), .IN2(n4304), .IN3(n4692), .Q(n4752) );
  NAND2X0 U9674 ( .IN1(g3167), .IN2(n1730), .QN(n3296) );
  NAND2X0 U9675 ( .IN1(g6565), .IN2(n5563), .QN(n3770) );
  NAND2X0 U9676 ( .IN1(g3873), .IN2(n5564), .QN(n3947) );
  NAND2X0 U9677 ( .IN1(g5873), .IN2(n5565), .QN(n3838) );
  NAND2X0 U9678 ( .IN1(g5527), .IN2(n5566), .QN(n3871) );
  NAND2X0 U9679 ( .IN1(g5180), .IN2(n5567), .QN(n3904) );
  NAND2X0 U9680 ( .IN1(g6219), .IN2(n5568), .QN(n3804) );
  NAND2X0 U9681 ( .IN1(g3522), .IN2(n5569), .QN(n3980) );
  NAND2X0 U9682 ( .IN1(g3171), .IN2(n5390), .QN(n4020) );
  NAND2X0 U9683 ( .IN1(g3530), .IN2(n5383), .QN(n3978) );
  NAND2X0 U9684 ( .IN1(g5188), .IN2(n5384), .QN(n3902) );
  NAND2X0 U9685 ( .IN1(g6227), .IN2(n5385), .QN(n3802) );
  NAND2X0 U9686 ( .IN1(g6573), .IN2(n5386), .QN(n3768) );
  NAND2X0 U9687 ( .IN1(g3881), .IN2(n5387), .QN(n3945) );
  NAND2X0 U9688 ( .IN1(test_so36), .IN2(n5388), .QN(n3836) );
  NAND2X0 U9689 ( .IN1(g5535), .IN2(n5389), .QN(n3869) );
  NOR2X0 U9690 ( .IN1(g25), .IN2(g22), .QN(g23190) );
  NAND2X0 U9691 ( .IN1(g3179), .IN2(g3171), .QN(n4017) );
  NAND2X0 U9692 ( .IN1(g5523), .IN2(n1968), .QN(n3289) );
  NAND2X0 U9693 ( .IN1(g5176), .IN2(n1581), .QN(n3287) );
  NAND2X0 U9694 ( .IN1(g6561), .IN2(n2224), .QN(n3295) );
  NAND2X0 U9695 ( .IN1(g3352), .IN2(n5400), .QN(n3089) );
  NAND2X0 U9696 ( .IN1(g6215), .IN2(n1514), .QN(n3292) );
  NAND2X0 U9697 ( .IN1(test_so33), .IN2(n1908), .QN(n3298) );
  NAND2X0 U9698 ( .IN1(g3518), .IN2(n1680), .QN(n3299) );
  NAND2X0 U9699 ( .IN1(g5869), .IN2(n1821), .QN(n3294) );
  OA21X1 U9700 ( .IN1(n4301), .IN2(n4692), .IN3(g4871), .Q(n3079) );
  OA21X1 U9701 ( .IN1(n4299), .IN2(n4692), .IN3(g4836), .Q(n3018) );
  OA21X1 U9702 ( .IN1(n4300), .IN2(n4692), .IN3(g4864), .Q(n3088) );
  OA21X1 U9703 ( .IN1(n4322), .IN2(n4698), .IN3(g4674), .Q(n3047) );
  OA21X1 U9704 ( .IN1(n4323), .IN2(n4698), .IN3(g4681), .Q(n3038) );
  NOR2X0 U9705 ( .IN1(n3711), .IN2(g5041), .QN(n3706) );
  NAND2X0 U9706 ( .IN1(g1183), .IN2(n5363), .QN(n3235) );
  OA21X1 U9707 ( .IN1(n5562), .IN2(g812), .IN3(g847), .Q(n4520) );
  NAND2X0 U9708 ( .IN1(g5357), .IN2(n5588), .QN(n3055) );
  NAND2X0 U9709 ( .IN1(test_so57), .IN2(n5589), .QN(n3037) );
  NAND2X0 U9710 ( .IN1(g6741), .IN2(n5590), .QN(n3017) );
  NAND2X0 U9711 ( .IN1(g3703), .IN2(n5591), .QN(n3078) );
  NAND2X0 U9712 ( .IN1(g6395), .IN2(n5592), .QN(n3028) );
  NAND2X0 U9713 ( .IN1(g5703), .IN2(n5593), .QN(n3046) );
  NAND2X0 U9714 ( .IN1(g4054), .IN2(n5594), .QN(n3070) );
  NAND2X0 U9715 ( .IN1(g3352), .IN2(g3288), .QN(n2741) );
  NAND2X0 U9716 ( .IN1(g6573), .IN2(g6565), .QN(n3776) );
  NAND2X0 U9717 ( .IN1(g5535), .IN2(g5527), .QN(n3877) );
  NAND2X0 U9718 ( .IN1(g5188), .IN2(g5180), .QN(n3910) );
  NAND2X0 U9719 ( .IN1(g3530), .IN2(g3522), .QN(n3986) );
  NAND2X0 U9720 ( .IN1(g3881), .IN2(g3873), .QN(n3953) );
  NAND2X0 U9721 ( .IN1(test_so36), .IN2(g5873), .QN(n3844) );
  NAND2X0 U9722 ( .IN1(g6227), .IN2(g6219), .QN(n3810) );
  OA21X1 U9723 ( .IN1(n3215), .IN2(n3216), .IN3(g17400), .Q(n3201) );
  NAND2X0 U9724 ( .IN1(test_so49), .IN2(n5364), .QN(n3155) );
  OA21X1 U9725 ( .IN1(n3235), .IN2(n3216), .IN3(g17316), .Q(n3221) );
  NAND2X0 U9726 ( .IN1(g691), .IN2(n5595), .QN(n2457) );
  OA21X1 U9727 ( .IN1(n3196), .IN2(g1171), .IN3(g1087), .Q(n3181) );
  NAND2X0 U9728 ( .IN1(g6741), .IN2(g6682), .QN(n2736) );
  NAND2X0 U9729 ( .IN1(g3703), .IN2(g3639), .QN(n2743) );
  NAND2X0 U9730 ( .IN1(g5703), .IN2(g5644), .QN(n2734) );
  NAND2X0 U9731 ( .IN1(g6395), .IN2(g6336), .QN(n2742) );
  NAND2X0 U9732 ( .IN1(g4785), .IN2(n5518), .QN(n2765) );
  NAND2X0 U9733 ( .IN1(g4975), .IN2(n5517), .QN(n2750) );
  NAND2X0 U9734 ( .IN1(n1609), .IN2(g4983), .QN(n2754) );
  NAND2X0 U9735 ( .IN1(n1728), .IN2(g4793), .QN(n2769) );
  NAND2X0 U9736 ( .IN1(test_so57), .IN2(g5990), .QN(n2745) );
  NAND2X0 U9737 ( .IN1(g5357), .IN2(g5297), .QN(n2739) );
  NAND2X0 U9738 ( .IN1(g4054), .IN2(g3990), .QN(n2746) );
  NAND2X0 U9739 ( .IN1(g13259), .IN2(n1696), .QN(n4492) );
  NAND2X0 U9740 ( .IN1(g13272), .IN2(n2034), .QN(n4468) );
  NAND2X0 U9741 ( .IN1(n1608), .IN2(g4966), .QN(n2751) );
  NAND2X0 U9742 ( .IN1(n1727), .IN2(g4776), .QN(n2766) );
  NAND2X0 U9743 ( .IN1(g1183), .IN2(g1171), .QN(n3215) );
  OR2X1 U9744 ( .IN1(n5380), .IN2(g4284), .Q(n4210) );
  NAND2X0 U9745 ( .IN1(g1668), .IN2(n5549), .QN(n2724) );
  NAND2X0 U9746 ( .IN1(g4087), .IN2(n5340), .QN(n3288) );
  NAND2X0 U9747 ( .IN1(g4093), .IN2(g4087), .QN(n3291) );
  NAND2X0 U9748 ( .IN1(g4093), .IN2(n5480), .QN(n3293) );
  OA22X1 U9749 ( .IN1(n4546), .IN2(n4547), .IN3(n4547), .IN4(n5358), .Q(n3676)
         );
  NOR2X0 U9750 ( .IN1(n4549), .IN2(n4548), .QN(n4546) );
  OA21X1 U9751 ( .IN1(n4548), .IN2(n4549), .IN3(g417), .Q(n4547) );
  AND3X1 U9752 ( .IN1(g392), .IN2(g405), .IN3(g401), .Q(n4549) );
  NOR2X0 U9753 ( .IN1(g24184), .IN2(n4881), .QN(n2417) );
  AND3X1 U9754 ( .IN1(n4882), .IN2(n4883), .IN3(n4884), .Q(n4881) );
  NAND4X0 U9755 ( .IN1(g4593), .IN2(g4584), .IN3(n5365), .IN4(n5274), .QN(
        n4883) );
  NAND3X0 U9756 ( .IN1(n5539), .IN2(n5303), .IN3(g4608), .QN(n4884) );
  OA21X1 U9757 ( .IN1(n3258), .IN2(g1367), .IN3(n3660), .Q(n3659) );
  OA21X1 U9758 ( .IN1(n3266), .IN2(g1024), .IN3(n3669), .Q(n3668) );
  NAND2X0 U9759 ( .IN1(g5041), .IN2(n1824), .QN(n3705) );
  NAND2X0 U9760 ( .IN1(g4709), .IN2(n5361), .QN(n2767) );
  NAND2X0 U9761 ( .IN1(g4899), .IN2(n5360), .QN(n2752) );
  NAND2X0 U9762 ( .IN1(n3472), .IN2(g4098), .QN(n3471) );
  NAND2X0 U9763 ( .IN1(test_so49), .IN2(g1514), .QN(n3135) );
  NAND2X0 U9764 ( .IN1(g2051), .IN2(n5371), .QN(n3599) );
  NAND2X0 U9765 ( .IN1(g2208), .IN2(n5376), .QN(n3580) );
  NAND2X0 U9766 ( .IN1(g2476), .IN2(n5373), .QN(n3542) );
  NAND2X0 U9767 ( .IN1(g1917), .IN2(n5374), .QN(n3617) );
  NAND2X0 U9768 ( .IN1(g2610), .IN2(n5372), .QN(n3523) );
  NAND2X0 U9769 ( .IN1(test_so21), .IN2(n5375), .QN(n3561) );
  NOR3X0 U9770 ( .IN1(n6002), .IN2(n6003), .IN3(n6004), .QN(g32185) );
  AO22X1 U9771 ( .IN1(g2927), .IN2(g2922), .IN3(g2941), .IN4(g2936), .Q(n6002)
         );
  AO22X1 U9772 ( .IN1(g2902), .IN2(test_so1), .IN3(g2917), .IN4(g2912), .Q(
        n6003) );
  AO222X1 U9773 ( .IN1(g2975), .IN2(g2970), .IN3(g2955), .IN4(g2950), .IN5(
        g2965), .IN6(test_so22), .Q(n6004) );
  NOR2X0 U9774 ( .IN1(n5359), .IN2(g1783), .QN(n3621) );
  NAND2X0 U9775 ( .IN1(test_so94), .IN2(n5370), .QN(n3652) );
  NAND2X0 U9776 ( .IN1(g3288), .IN2(n5604), .QN(n3090) );
  NAND2X0 U9777 ( .IN1(g5297), .IN2(n5393), .QN(n3056) );
  NAND2X0 U9778 ( .IN1(g5990), .IN2(n5394), .QN(n3039) );
  NAND2X0 U9779 ( .IN1(g3990), .IN2(n5395), .QN(n3071) );
  NAND2X0 U9780 ( .IN1(g6336), .IN2(n5396), .QN(n3029) );
  NAND2X0 U9781 ( .IN1(g5644), .IN2(n5397), .QN(n3048) );
  NAND2X0 U9782 ( .IN1(g6682), .IN2(n5398), .QN(n3019) );
  NAND2X0 U9783 ( .IN1(g3639), .IN2(n5399), .QN(n3080) );
  NAND2X0 U9784 ( .IN1(g4064), .IN2(g4057), .QN(n4723) );
  NAND2X0 U9785 ( .IN1(g703), .IN2(n4531), .QN(n4527) );
  NAND4X0 U9786 ( .IN1(g681), .IN2(n4532), .IN3(test_so87), .IN4(n4533), .QN(
        n4531) );
  NOR4X0 U9787 ( .IN1(g650), .IN2(g645), .IN3(n4534), .IN4(n4535), .QN(n4533)
         );
  NAND2X0 U9788 ( .IN1(g5046), .IN2(n1823), .QN(n3697) );
  NAND2X0 U9789 ( .IN1(test_so94), .IN2(n5525), .QN(n3004) );
  NAND3X0 U9790 ( .IN1(n5363), .IN2(n5599), .IN3(g13259), .QN(n4499) );
  NAND3X0 U9791 ( .IN1(DFF_178_n1), .IN2(n5636), .IN3(n2668), .QN(n2675) );
  NAND3X0 U9792 ( .IN1(DFF_672_n1), .IN2(n5637), .IN3(n2668), .QN(n2654) );
  NAND2X0 U9793 ( .IN1(g1270), .IN2(n3662), .QN(n3262) );
  NAND2X0 U9794 ( .IN1(g925), .IN2(n3671), .QN(n3270) );
  OA21X1 U9795 ( .IN1(n3135), .IN2(n3136), .IN3(g17423), .Q(n3122) );
  AO21X1 U9796 ( .IN1(g4616), .IN2(n2601), .IN3(n1299), .Q(n2592) );
  NAND2X0 U9797 ( .IN1(g4082), .IN2(n4729), .QN(n4328) );
  NAND2X0 U9798 ( .IN1(n2583), .IN2(g4340), .QN(n2693) );
  NAND2X0 U9799 ( .IN1(n3942), .IN2(g4087), .QN(n3729) );
  NAND2X0 U9800 ( .IN1(g2729), .IN2(g2724), .QN(n2632) );
  NOR2X0 U9801 ( .IN1(n5508), .IN2(g2610), .QN(n3510) );
  OA21X1 U9802 ( .IN1(n3155), .IN2(n3136), .IN3(g17404), .Q(n3141) );
  OA21X1 U9803 ( .IN1(n5364), .IN2(n3117), .IN3(g17320), .Q(n3160) );
  NOR2X0 U9804 ( .IN1(n5507), .IN2(g2051), .QN(n3585) );
  NOR2X0 U9805 ( .IN1(n5509), .IN2(g2476), .QN(n3529) );
  NOR2X0 U9806 ( .IN1(n5510), .IN2(g1917), .QN(n3603) );
  NOR2X0 U9807 ( .IN1(n5511), .IN2(test_so21), .QN(n3547) );
  NOR2X0 U9808 ( .IN1(n5512), .IN2(g2208), .QN(n3566) );
  NAND4X0 U9809 ( .IN1(n5412), .IN2(n5626), .IN3(n4982), .IN4(n4983), .QN(
        n2440) );
  NOR2X0 U9810 ( .IN1(g1858), .IN2(g1844), .QN(n4982) );
  NOR4X0 U9811 ( .IN1(g2126), .IN2(g2112), .IN3(g1992), .IN4(g1978), .QN(n4983) );
  OA21X1 U9812 ( .IN1(n3117), .IN2(g1514), .IN3(g1430), .Q(n3102) );
  NAND3X0 U9813 ( .IN1(n2760), .IN2(n2761), .IN3(g63), .QN(n2669) );
  NAND3X0 U9814 ( .IN1(n2760), .IN2(n2775), .IN3(g63), .QN(n2689) );
  NAND4X0 U9815 ( .IN1(n5621), .IN2(n5407), .IN3(n4978), .IN4(n4979), .QN(
        n2433) );
  NOR2X0 U9816 ( .IN1(g1798), .IN2(g1779), .QN(n4978) );
  NOR4X0 U9817 ( .IN1(g2066), .IN2(g2047), .IN3(g1932), .IN4(g1913), .QN(n4979) );
  NOR2X0 U9818 ( .IN1(n5525), .IN2(test_so94), .QN(n3639) );
  NOR2X0 U9819 ( .IN1(n3698), .IN2(g5052), .QN(n3452) );
  AO221X1 U9820 ( .IN1(n4822), .IN2(n5520), .IN3(g691), .IN4(n4823), .IN5(
        n4824), .Q(n4821) );
  NAND2X0 U9821 ( .IN1(n5481), .IN2(n5287), .QN(n4823) );
  OR3X1 U9822 ( .IN1(g411), .IN2(g424), .IN3(n5358), .Q(n4822) );
  NAND3X0 U9823 ( .IN1(n5364), .IN2(n5542), .IN3(g13272), .QN(n4475) );
  NOR2X0 U9824 ( .IN1(g4082), .IN2(g4141), .QN(n4724) );
  ISOLANDX1 U9825 ( .D(g112), .ISO(n1300), .Q(n3115) );
  AND3X1 U9826 ( .IN1(g904), .IN2(g12919), .IN3(g921), .Q(n4811) );
  NAND3X0 U9827 ( .IN1(n1499), .IN2(g1657), .IN3(g1624), .QN(n4151) );
  NAND3X0 U9828 ( .IN1(n1713), .IN2(g2619), .IN3(g2587), .QN(n4067) );
  NAND3X0 U9829 ( .IN1(n1863), .IN2(g2217), .IN3(g2185), .QN(n4103) );
  NAND3X0 U9830 ( .IN1(n1770), .IN2(g1926), .IN3(g1894), .QN(n4127) );
  NAND3X0 U9831 ( .IN1(n1859), .IN2(g2060), .IN3(g2028), .QN(n4115) );
  NAND3X0 U9832 ( .IN1(n1762), .IN2(g2485), .IN3(g2453), .QN(n4079) );
  AND3X1 U9833 ( .IN1(g1266), .IN2(g1249), .IN3(g12923), .Q(n4804) );
  NOR2X0 U9834 ( .IN1(g3143), .IN2(g3129), .QN(n2469) );
  NAND3X0 U9835 ( .IN1(n2668), .IN2(n5541), .IN3(g4507), .QN(g33874) );
  AND3X1 U9836 ( .IN1(g12919), .IN2(n5084), .IN3(g1052), .Q(n4936) );
  AND3X1 U9837 ( .IN1(g12923), .IN2(n5060), .IN3(g1395), .Q(n4911) );
  AND3X1 U9838 ( .IN1(n5368), .IN2(n5285), .IN3(g4776), .Q(n4317) );
  AND3X1 U9839 ( .IN1(n5367), .IN2(n5284), .IN3(g4966), .Q(n4295) );
  NAND3X0 U9840 ( .IN1(g1171), .IN2(n5599), .IN3(g13259), .QN(n4509) );
  NAND3X0 U9841 ( .IN1(g1514), .IN2(n5542), .IN3(g13272), .QN(n4485) );
  AO22X1 U9842 ( .IN1(g437), .IN2(n4550), .IN3(n4551), .IN4(g424), .Q(n4548)
         );
  NOR2X0 U9843 ( .IN1(g405), .IN2(g392), .QN(n4551) );
  XOR2X1 U9844 ( .IN1(g405), .IN2(g392), .Q(n4550) );
  NOR2X0 U9845 ( .IN1(g3167), .IN2(n1280), .QN(n3494) );
  AND3X1 U9846 ( .IN1(g5041), .IN2(g24168), .IN3(n4672), .Q(n3721) );
  NOR2X0 U9847 ( .IN1(n3693), .IN2(g5033), .QN(n3688) );
  NAND2X0 U9848 ( .IN1(n3282), .IN2(n3283), .QN(n2515) );
  OAI22X1 U9849 ( .IN1(n3284), .IN2(n5350), .IN3(g4098), .IN4(n3285), .QN(
        n3283) );
  OA221X1 U9850 ( .IN1(n3286), .IN2(n3287), .IN3(n3288), .IN4(n3289), .IN5(
        n3290), .Q(n3285) );
  OA221X1 U9851 ( .IN1(n3286), .IN2(n3295), .IN3(n3288), .IN4(n3296), .IN5(
        n3297), .Q(n3284) );
  AND3X1 U9852 ( .IN1(g385), .IN2(g376), .IN3(g8719), .Q(n2642) );
  NAND3X0 U9853 ( .IN1(g518), .IN2(n5548), .IN3(g203), .QN(n4203) );
  AND3X1 U9854 ( .IN1(g5052), .IN2(n5950), .IN3(n4672), .Q(n3722) );
  NAND3X0 U9855 ( .IN1(g5029), .IN2(g5016), .IN3(g5062), .QN(n3692) );
  NAND3X0 U9856 ( .IN1(g2729), .IN2(g2735), .IN3(n4064), .QN(n3506) );
  NAND3X0 U9857 ( .IN1(g518), .IN2(n5548), .IN3(n2075), .QN(n4829) );
  NAND2X0 U9858 ( .IN1(g112), .IN2(g31862), .QN(n3240) );
  NAND4X0 U9859 ( .IN1(g12238), .IN2(g17519), .IN3(g17674), .IN4(g14662), .QN(
        n5160) );
  NAND4X0 U9860 ( .IN1(g12300), .IN2(g17580), .IN3(g17711), .IN4(g14694), .QN(
        n5155) );
  NAND4X0 U9861 ( .IN1(g12470), .IN2(g17688), .IN3(g17778), .IN4(g14828), .QN(
        n5140) );
  NAND4X0 U9862 ( .IN1(g12350), .IN2(g17607), .IN3(g17739), .IN4(g14738), .QN(
        n5150) );
  NAND4X0 U9863 ( .IN1(g11418), .IN2(g16659), .IN3(g16775), .IN4(g13966), .QN(
        n5182) );
  NAND4X0 U9864 ( .IN1(g12422), .IN2(g17649), .IN3(g17760), .IN4(g14779), .QN(
        n5145) );
  NAND4X0 U9865 ( .IN1(g11349), .IN2(g16603), .IN3(g16718), .IN4(g13895), .QN(
        n5192) );
  NAND4X0 U9866 ( .IN1(g11388), .IN2(g16627), .IN3(g16744), .IN4(g13926), .QN(
        n5187) );
  NAND2X0 U9867 ( .IN1(g1300), .IN2(n4475), .QN(n5056) );
  OA21X1 U9868 ( .IN1(n3258), .IN2(g1345), .IN3(n4176), .Q(n3734) );
  OA21X1 U9869 ( .IN1(n3266), .IN2(g1002), .IN3(n4194), .Q(n3739) );
  OA21X1 U9870 ( .IN1(n3258), .IN2(g1361), .IN3(n3734), .Q(n3660) );
  OA21X1 U9871 ( .IN1(n3266), .IN2(g1018), .IN3(n3739), .Q(n3669) );
  NAND3X0 U9872 ( .IN1(n3505), .IN2(test_so30), .IN3(g2735), .QN(n2631) );
  AND3X1 U9873 ( .IN1(g817), .IN2(n4948), .IN3(g832), .Q(n4814) );
  NAND4X0 U9874 ( .IN1(g262), .IN2(g255), .IN3(g269), .IN4(n5128), .QN(n4834)
         );
  NOR4X0 U9875 ( .IN1(g246), .IN2(g239), .IN3(g232), .IN4(g225), .QN(n5128) );
  NAND3X0 U9876 ( .IN1(g5033), .IN2(n1874), .IN3(g5037), .QN(n3710) );
  NAND3X0 U9877 ( .IN1(g2051), .IN2(n5507), .IN3(n1859), .QN(n4123) );
  NAND3X0 U9878 ( .IN1(g2610), .IN2(n5508), .IN3(n1713), .QN(n4075) );
  NAND3X0 U9879 ( .IN1(g2476), .IN2(n5509), .IN3(n1762), .QN(n4087) );
  NAND3X0 U9880 ( .IN1(g1917), .IN2(n5510), .IN3(n1770), .QN(n4135) );
  NAND3X0 U9881 ( .IN1(g2208), .IN2(n5512), .IN3(n1863), .QN(n4111) );
  NAND4X0 U9882 ( .IN1(test_so68), .IN2(n5546), .IN3(g1404), .IN4(n3175), .QN(
        n3136) );
  NOR3X0 U9883 ( .IN1(g1554), .IN2(g1564), .IN3(g1559), .QN(n3175) );
  NAND4X0 U9884 ( .IN1(g1061), .IN2(n5547), .IN3(g979), .IN4(n5264), .QN(n3216) );
  NOR3X0 U9885 ( .IN1(test_so76), .IN2(g1221), .IN3(g1216), .QN(n5264) );
  ISOLANDX1 U9886 ( .D(g370), .ISO(n5121), .Q(n4948) );
  AO221X1 U9887 ( .IN1(n4775), .IN2(n4776), .IN3(n1946), .IN4(n4777), .IN5(
        n4778), .Q(n4373) );
  INVX0 U9888 ( .IN(n4775), .QN(n1946) );
  XNOR2X1 U9889 ( .IN1(g11349), .IN2(n5527), .Q(n4775) );
  NAND3X0 U9890 ( .IN1(n4791), .IN2(n4792), .IN3(n4793), .QN(n4777) );
  AO221X1 U9891 ( .IN1(n4646), .IN2(n4647), .IN3(n1635), .IN4(n4648), .IN5(
        n4649), .Q(n4282) );
  NAND3X0 U9892 ( .IN1(n4663), .IN2(n4664), .IN3(n4665), .QN(n4648) );
  INVX0 U9893 ( .IN(n4646), .QN(n1635) );
  XNOR2X1 U9894 ( .IN1(g12238), .IN2(n5515), .Q(n4646) );
  AO221X1 U9895 ( .IN1(n4600), .IN2(n4601), .IN3(n1522), .IN4(n4602), .IN5(
        n4603), .Q(n4252) );
  INVX0 U9896 ( .IN(n4600), .QN(n1522) );
  XNOR2X1 U9897 ( .IN1(g12350), .IN2(n5528), .Q(n4600) );
  NAND3X0 U9898 ( .IN1(n4617), .IN2(n4618), .IN3(n4619), .QN(n4602) );
  AO221X1 U9899 ( .IN1(n4623), .IN2(n4624), .IN3(n1534), .IN4(n4625), .IN5(
        n4626), .Q(n4267) );
  INVX0 U9900 ( .IN(n4623), .QN(n1534) );
  XNOR2X1 U9901 ( .IN1(g12300), .IN2(n5529), .Q(n4623) );
  NAND3X0 U9902 ( .IN1(n4640), .IN2(n4641), .IN3(n4642), .QN(n4625) );
  AO221X1 U9903 ( .IN1(n4730), .IN2(n4731), .IN3(n1504), .IN4(n4732), .IN5(
        n4733), .Q(n4343) );
  INVX0 U9904 ( .IN(n4730), .QN(n1504) );
  XNOR2X1 U9905 ( .IN1(g11418), .IN2(n5530), .Q(n4730) );
  NAND3X0 U9906 ( .IN1(n4746), .IN2(n4747), .IN3(n4748), .QN(n4732) );
  AO221X1 U9907 ( .IN1(n4554), .IN2(n4555), .IN3(n1676), .IN4(n4556), .IN5(
        n4557), .Q(n4222) );
  INVX0 U9908 ( .IN(n4554), .QN(n1676) );
  XNOR2X1 U9909 ( .IN1(g12470), .IN2(n5531), .Q(n4554) );
  NAND3X0 U9910 ( .IN1(n4571), .IN2(n4572), .IN3(n4573), .QN(n4556) );
  AO221X1 U9911 ( .IN1(n4753), .IN2(n4754), .IN3(n2011), .IN4(n4755), .IN5(
        n4756), .Q(n4358) );
  INVX0 U9912 ( .IN(n4753), .QN(n2011) );
  XNOR2X1 U9913 ( .IN1(g11388), .IN2(n5532), .Q(n4753) );
  NAND3X0 U9914 ( .IN1(n4769), .IN2(n4770), .IN3(n4771), .QN(n4755) );
  AO221X1 U9915 ( .IN1(n4577), .IN2(n4578), .IN3(n1954), .IN4(n4579), .IN5(
        n4580), .Q(n4237) );
  INVX0 U9916 ( .IN(n4577), .QN(n1954) );
  XNOR2X1 U9917 ( .IN1(g12422), .IN2(n5533), .Q(n4577) );
  NAND3X0 U9918 ( .IN1(n4594), .IN2(n4595), .IN3(n4596), .QN(n4579) );
  AND3X1 U9919 ( .IN1(n2760), .IN2(n3282), .IN3(g43), .Q(n3933) );
  NAND2X0 U9920 ( .IN1(g2729), .IN2(n5301), .QN(n2637) );
  AND3X1 U9921 ( .IN1(g5062), .IN2(n5615), .IN3(g5046), .Q(n4672) );
  AND3X1 U9922 ( .IN1(g996), .IN2(n5642), .IN3(g1178), .Q(n4919) );
  AO22X1 U9923 ( .IN1(g24179), .IN2(g4146), .IN3(g24178), .IN4(n5981), .Q(
        n3939) );
  AO22X1 U9924 ( .IN1(g24177), .IN2(g4157), .IN3(g24175), .IN4(n5983), .Q(
        n3938) );
  AND3X1 U9925 ( .IN1(g5022), .IN2(n5578), .IN3(g5057), .Q(n4670) );
  NAND2X0 U9926 ( .IN1(n2790), .IN2(test_so30), .QN(n2789) );
  ISOLANDX1 U9927 ( .D(n3933), .ISO(g4098), .Q(n3833) );
  NOR2X0 U9928 ( .IN1(n6005), .IN2(n1300), .QN(n2613) );
  NOR2X0 U9929 ( .IN1(n6006), .IN2(n1300), .QN(n2629) );
  OR2X1 U9930 ( .IN1(n5571), .IN2(g6555), .Q(n3407) );
  OR2X1 U9931 ( .IN1(n5572), .IN2(g3863), .Q(n3482) );
  OR2X1 U9932 ( .IN1(n5573), .IN2(g5863), .Q(n3427) );
  OR2X1 U9933 ( .IN1(n5575), .IN2(g5517), .Q(n3437) );
  OR2X1 U9934 ( .IN1(n5574), .IN2(g6209), .Q(n3417) );
  OR2X1 U9935 ( .IN1(n5576), .IN2(g3512), .Q(n3492) );
  OR2X1 U9936 ( .IN1(n5570), .IN2(g5170), .Q(n3447) );
  NOR2X0 U9937 ( .IN1(g1373), .IN2(n3258), .QN(n3257) );
  NOR2X0 U9938 ( .IN1(g1030), .IN2(n3266), .QN(n3265) );
  AO221X1 U9939 ( .IN1(g1677), .IN2(n5299), .IN3(g1811), .IN4(g2715), .IN5(
        g2719), .Q(n4059) );
  AO221X1 U9940 ( .IN1(g2236), .IN2(n5299), .IN3(g2370), .IN4(g2715), .IN5(
        g2719), .Q(n4047) );
  NAND3X0 U9941 ( .IN1(g4322), .IN2(g4332), .IN3(n2607), .QN(n2604) );
  NAND2X0 U9942 ( .IN1(g1389), .IN2(n5067), .QN(n4800) );
  XNOR2X1 U9943 ( .IN1(g191), .IN2(g8358), .Q(n5130) );
  NAND2X0 U9944 ( .IN1(g1373), .IN2(g1361), .QN(n5066) );
  NAND2X0 U9945 ( .IN1(g1030), .IN2(g1018), .QN(n5090) );
  NAND4X0 U9946 ( .IN1(DFF_1234_n1), .IN2(DFF_909_n1), .IN3(DFF_480_n1), .IN4(
        n5256), .QN(n5255) );
  NOR4X0 U9947 ( .IN1(g8789), .IN2(g8788), .IN3(g8787), .IN4(g8785), .QN(n5256) );
  NAND3X0 U9948 ( .IN1(g17577), .IN2(g31860), .IN3(g25219), .QN(n4279) );
  NAND2X0 U9949 ( .IN1(g4944), .IN2(n2135), .QN(n4301) );
  NAND2X0 U9950 ( .IN1(g4754), .IN2(n2101), .QN(n4323) );
  NAND2X0 U9951 ( .IN1(g4933), .IN2(n2136), .QN(n4300) );
  NAND2X0 U9952 ( .IN1(g4743), .IN2(n2103), .QN(n4322) );
  ISOLANDX1 U9953 ( .D(g671), .ISO(n1538), .Q(n4526) );
  OA22X1 U9954 ( .IN1(g4512), .IN2(g4581), .IN3(n3062), .IN4(n5670), .Q(n2779)
         );
  OR2X1 U9955 ( .IN1(g20049), .IN2(n2416), .Q(n3062) );
  NOR2X0 U9956 ( .IN1(n6007), .IN2(g4427), .QN(n2479) );
  ISOLANDX1 U9957 ( .D(g4843), .ISO(n5283), .Q(n2563) );
  ISOLANDX1 U9958 ( .D(test_so19), .ISO(n5656), .Q(n2573) );
  OA22X1 U9959 ( .IN1(g4552), .IN2(g4581), .IN3(n3061), .IN4(n5670), .Q(n2784)
         );
  OR2X1 U9960 ( .IN1(g4575), .IN2(n2416), .Q(n3061) );
  NAND3X0 U9961 ( .IN1(g17604), .IN2(n2307), .IN3(g5689), .QN(n4264) );
  NAND3X0 U9962 ( .IN1(g16624), .IN2(n1880), .IN3(g3338), .QN(n4370) );
  NAND3X0 U9963 ( .IN1(g17722), .IN2(n2123), .IN3(g6727), .QN(n4219) );
  NAND3X0 U9964 ( .IN1(g16693), .IN2(n1747), .IN3(g4040), .QN(n4340) );
  NAND3X0 U9965 ( .IN1(g17646), .IN2(n1870), .IN3(g6035), .QN(n4249) );
  NAND3X0 U9966 ( .IN1(g16656), .IN2(n1940), .IN3(g3689), .QN(n4355) );
  NAND3X0 U9967 ( .IN1(g17685), .IN2(n1625), .IN3(test_so69), .QN(n4234) );
  ISOLANDX1 U9968 ( .D(n3084), .ISO(g4358), .Q(n3023) );
  NAND3X0 U9969 ( .IN1(g482), .IN2(n5327), .IN3(g490), .QN(n4828) );
  NAND4X0 U9970 ( .IN1(g703), .IN2(test_so87), .IN3(n5112), .IN4(n5113), .QN(
        n4819) );
  NOR4X0 U9971 ( .IN1(g691), .IN2(g650), .IN3(g645), .IN4(n4534), .QN(n5113)
         );
  ISOLANDX1 U9972 ( .D(g681), .ISO(n4535), .Q(n5112) );
  NOR3X0 U9973 ( .IN1(g3161), .IN2(g3167), .IN3(g3155), .QN(n4034) );
  NOR3X0 U9974 ( .IN1(g6555), .IN2(g6561), .IN3(g6549), .QN(n3792) );
  NOR3X0 U9975 ( .IN1(g5170), .IN2(g5176), .IN3(g5164), .QN(n3926) );
  NOR3X0 U9976 ( .IN1(g6209), .IN2(g6215), .IN3(g6203), .QN(n3826) );
  NOR3X0 U9977 ( .IN1(g5517), .IN2(g5523), .IN3(g5511), .QN(n3893) );
  NOR3X0 U9978 ( .IN1(g3863), .IN2(test_so33), .IN3(g3857), .QN(n3969) );
  NOR3X0 U9979 ( .IN1(g5863), .IN2(g5869), .IN3(g5857), .QN(n3860) );
  NOR3X0 U9980 ( .IN1(g3512), .IN2(g3518), .IN3(g3506), .QN(n4002) );
  AND2X1 U9981 ( .IN1(g1542), .IN2(n4166), .Q(n4163) );
  AND2X1 U9982 ( .IN1(g1199), .IN2(n4184), .Q(n4181) );
  XOR3X1 U9983 ( .IN1(g255), .IN2(n6008), .IN3(n6009), .Q(n5106) );
  XNOR2X1 U9984 ( .IN1(g269), .IN2(g262), .Q(n6009) );
  OR3X1 U9985 ( .IN1(n4492), .IN2(g1105), .IN3(n4924), .Q(n4933) );
  NOR2X0 U9986 ( .IN1(n6010), .IN2(n1300), .QN(n3084) );
  NAND3X0 U9987 ( .IN1(g1936), .IN2(n5503), .IN3(g112), .QN(n3202) );
  NAND3X0 U9988 ( .IN1(g2361), .IN2(n5513), .IN3(g112), .QN(n3142) );
  NAND3X0 U9989 ( .IN1(g2227), .IN2(n5514), .IN3(g112), .QN(n3161) );
  NAND3X0 U9990 ( .IN1(g1802), .IN2(n5504), .IN3(g112), .QN(n3222) );
  NAND3X0 U9991 ( .IN1(g2070), .IN2(n5505), .IN3(g112), .QN(n3182) );
  ISOLANDX1 U9992 ( .D(n3675), .ISO(n3676), .Q(n2644) );
  NAND4X0 U9993 ( .IN1(n3677), .IN2(n3678), .IN3(n5358), .IN4(n5520), .QN(
        n3675) );
  OAI21X1 U9994 ( .IN1(n3680), .IN2(g441), .IN3(g392), .QN(n3677) );
  AO21X1 U9995 ( .IN1(n3679), .IN2(n5629), .IN3(g392), .Q(n3678) );
  NAND3X0 U9996 ( .IN1(g2495), .IN2(n5523), .IN3(g112), .QN(n3123) );
  NAND3X0 U9997 ( .IN1(g2629), .IN2(n5524), .IN3(g112), .QN(n3103) );
  OR3X1 U9998 ( .IN1(n4475), .IN2(g1300), .IN3(n4899), .Q(n5058) );
  OR3X1 U9999 ( .IN1(n4468), .IN2(g1448), .IN3(n4899), .Q(n4908) );
  NOR3X0 U10000 ( .IN1(n5301), .IN2(g2729), .IN3(n2631), .QN(n2618) );
  NAND4X0 U10001 ( .IN1(g239), .IN2(g232), .IN3(g246), .IN4(n5127), .QN(n4835)
         );
  NOR4X0 U10002 ( .IN1(g269), .IN2(g262), .IN3(g255), .IN4(n5597), .QN(n5127)
         );
  NAND3X0 U10003 ( .IN1(n5369), .IN2(n5601), .IN3(g5022), .QN(n3693) );
  NOR2X0 U10004 ( .IN1(n4542), .IN2(n5820), .QN(n4538) );
  NAND3X0 U10005 ( .IN1(g358), .IN2(n5633), .IN3(g385), .QN(n4818) );
  NAND4X0 U10006 ( .IN1(g370), .IN2(g8719), .IN3(g376), .IN4(n5632), .QN(n2645) );
  NAND3X0 U10007 ( .IN1(n2702), .IN2(n5849), .IN3(g26960), .QN(n2697) );
  AO21X1 U10008 ( .IN1(n2668), .IN2(n5846), .IN3(n2416), .Q(n2702) );
  XOR2X1 U10009 ( .IN1(g728), .IN2(g661), .Q(n4534) );
  OA22X1 U10010 ( .IN1(n4789), .IN2(n3089), .IN3(n4790), .IN4(n2741), .Q(n4788) );
  AOI22X1 U10011 ( .IN1(g3247), .IN2(g16686), .IN3(g3263), .IN4(g16624), .QN(
        n4790) );
  AOI22X1 U10012 ( .IN1(g3191), .IN2(g11349), .IN3(g3215), .IN4(g16874), .QN(
        n4789) );
  OA22X1 U10013 ( .IN1(n4638), .IN2(n3046), .IN3(n4639), .IN4(n2734), .Q(n4637) );
  AOI22X1 U10014 ( .IN1(g5603), .IN2(g17678), .IN3(g5619), .IN4(g17604), .QN(
        n4639) );
  AOI22X1 U10015 ( .IN1(g5547), .IN2(g12300), .IN3(g5571), .IN4(g17813), .QN(
        n4638) );
  OA22X1 U10016 ( .IN1(n4569), .IN2(n3017), .IN3(n4570), .IN4(n2736), .Q(n4568) );
  AOI22X1 U10017 ( .IN1(g6641), .IN2(g17764), .IN3(g6657), .IN4(g17722), .QN(
        n4570) );
  AOI22X1 U10018 ( .IN1(test_so71), .IN2(g12470), .IN3(g6609), .IN4(g17871), 
        .QN(n4569) );
  OA22X1 U10019 ( .IN1(n4767), .IN2(n3078), .IN3(n4768), .IN4(n2743), .Q(n4766) );
  AOI22X1 U10020 ( .IN1(g3598), .IN2(g16722), .IN3(g3614), .IN4(g16656), .QN(
        n4768) );
  AOI22X1 U10021 ( .IN1(g3542), .IN2(g11388), .IN3(g3566), .IN4(g16924), .QN(
        n4767) );
  OA22X1 U10022 ( .IN1(n4592), .IN2(n3028), .IN3(n4593), .IN4(n2742), .Q(n4591) );
  AOI22X1 U10023 ( .IN1(g6295), .IN2(g17743), .IN3(g6311), .IN4(g17685), .QN(
        n4593) );
  AOI22X1 U10024 ( .IN1(g6239), .IN2(g12422), .IN3(g6263), .IN4(g17845), .QN(
        n4592) );
  OA22X1 U10025 ( .IN1(n4661), .IN2(n3055), .IN3(n4662), .IN4(n2739), .Q(n4660) );
  AOI22X1 U10026 ( .IN1(g5256), .IN2(g17639), .IN3(g5272), .IN4(g17577), .QN(
        n4662) );
  AOI22X1 U10027 ( .IN1(g5200), .IN2(g12238), .IN3(g5224), .IN4(g17787), .QN(
        n4661) );
  OA22X1 U10028 ( .IN1(n4615), .IN2(n3037), .IN3(n4616), .IN4(n2745), .Q(n4614) );
  AOI22X1 U10029 ( .IN1(g5949), .IN2(g17715), .IN3(test_so13), .IN4(g17646), 
        .QN(n4616) );
  AOI22X1 U10030 ( .IN1(g5893), .IN2(g12350), .IN3(test_so28), .IN4(g17819), 
        .QN(n4615) );
  OA22X1 U10031 ( .IN1(n4744), .IN2(n3070), .IN3(n4745), .IN4(n2746), .Q(n4743) );
  AOI22X1 U10032 ( .IN1(test_so65), .IN2(g16748), .IN3(g3965), .IN4(g16693), 
        .QN(n4745) );
  AOI22X1 U10033 ( .IN1(g3893), .IN2(g11418), .IN3(g3917), .IN4(g16955), .QN(
        n4744) );
  XOR2X1 U10034 ( .IN1(g655), .IN2(g718), .Q(n4535) );
  NOR3X0 U10035 ( .IN1(n5391), .IN2(g4639), .IN3(n5309), .QN(n2583) );
  NAND3X0 U10036 ( .IN1(g2236), .IN2(n3580), .IN3(g2250), .QN(n4415) );
  NAND3X0 U10037 ( .IN1(g1811), .IN2(n3634), .IN3(g1825), .QN(n4448) );
  NAND3X0 U10038 ( .IN1(g2370), .IN2(n3561), .IN3(g2384), .QN(n4403) );
  NAND3X0 U10039 ( .IN1(g1677), .IN2(n3652), .IN3(g1691), .QN(n4459) );
  NAND3X0 U10040 ( .IN1(test_so78), .IN2(n3599), .IN3(g2079), .QN(n4426) );
  NAND3X0 U10041 ( .IN1(g1959), .IN2(n3617), .IN3(test_so53), .QN(n4437) );
  NAND3X0 U10042 ( .IN1(g2518), .IN2(n3542), .IN3(g2504), .QN(n4392) );
  NAND3X0 U10043 ( .IN1(g2652), .IN2(n3523), .IN3(g2638), .QN(n4380) );
  NAND3X0 U10044 ( .IN1(n5517), .IN2(n5360), .IN3(g4888), .QN(n4299) );
  NAND3X0 U10045 ( .IN1(n5518), .IN2(n5361), .IN3(g4698), .QN(n4321) );
  NAND3X0 U10046 ( .IN1(g4639), .IN2(n1298), .IN3(test_so3), .QN(n2586) );
  OR2X1 U10047 ( .IN1(n3216), .IN2(g1183), .Q(n3196) );
  NOR2X0 U10048 ( .IN1(n5178), .IN2(g4235), .QN(n5177) );
  NOR4X0 U10049 ( .IN1(n5179), .IN2(g11770), .IN3(g8916), .IN4(g8915), .QN(
        n5178) );
  NAND4X0 U10050 ( .IN1(DFF_992_n1), .IN2(DFF_418_n1), .IN3(DFF_944_n1), .IN4(
        DFF_1338_n1), .QN(n5179) );
  OR2X1 U10051 ( .IN1(n3136), .IN2(test_so49), .Q(n3117) );
  NAND2X0 U10052 ( .IN1(g101), .IN2(n1381), .QN(n2674) );
  NAND2X0 U10053 ( .IN1(g71), .IN2(n1386), .QN(n2653) );
  NAND3X0 U10054 ( .IN1(g13895), .IN2(g3219), .IN3(n1881), .QN(n4791) );
  NAND3X0 U10055 ( .IN1(g14662), .IN2(test_so82), .IN3(n1893), .QN(n4663) );
  NAND3X0 U10056 ( .IN1(g14738), .IN2(g5921), .IN3(n1869), .QN(n4617) );
  NAND3X0 U10057 ( .IN1(g14694), .IN2(g5575), .IN3(n2304), .QN(n4640) );
  NAND3X0 U10058 ( .IN1(g13966), .IN2(g3921), .IN3(n1749), .QN(n4746) );
  NAND3X0 U10059 ( .IN1(g14828), .IN2(g6613), .IN3(n2122), .QN(n4571) );
  NAND3X0 U10060 ( .IN1(g13926), .IN2(g3570), .IN3(n1941), .QN(n4769) );
  NAND3X0 U10061 ( .IN1(g14779), .IN2(g6267), .IN3(n1624), .QN(n4594) );
  NAND3X0 U10062 ( .IN1(n4794), .IN2(n4795), .IN3(n4796), .QN(n4776) );
  NAND3X0 U10063 ( .IN1(n1881), .IN2(test_so84), .IN3(g16603), .QN(n4796) );
  NAND3X0 U10064 ( .IN1(g3243), .IN2(n1882), .IN3(g16718), .QN(n4794) );
  NAND3X0 U10065 ( .IN1(n1883), .IN2(g3227), .IN3(g13895), .QN(n4795) );
  NAND3X0 U10066 ( .IN1(n4666), .IN2(n4667), .IN3(n4668), .QN(n4647) );
  NAND3X0 U10067 ( .IN1(n1893), .IN2(g5268), .IN3(g17519), .QN(n4668) );
  NAND3X0 U10068 ( .IN1(g5252), .IN2(n1891), .IN3(g17674), .QN(n4666) );
  NAND3X0 U10069 ( .IN1(n1890), .IN2(g5236), .IN3(g14662), .QN(n4667) );
  NAND3X0 U10070 ( .IN1(n4620), .IN2(n4621), .IN3(n4622), .QN(n4601) );
  NAND3X0 U10071 ( .IN1(n1869), .IN2(g5961), .IN3(g17607), .QN(n4622) );
  NAND3X0 U10072 ( .IN1(g5945), .IN2(n1867), .IN3(g17739), .QN(n4620) );
  NAND3X0 U10073 ( .IN1(n1866), .IN2(g5929), .IN3(g14738), .QN(n4621) );
  NAND3X0 U10074 ( .IN1(n4643), .IN2(n4644), .IN3(n4645), .QN(n4624) );
  NAND3X0 U10075 ( .IN1(n2304), .IN2(g5615), .IN3(g17580), .QN(n4645) );
  NAND3X0 U10076 ( .IN1(g5599), .IN2(n2303), .IN3(g17711), .QN(n4643) );
  NAND3X0 U10077 ( .IN1(n2305), .IN2(g5583), .IN3(g14694), .QN(n4644) );
  NAND3X0 U10078 ( .IN1(n4749), .IN2(n4750), .IN3(n4751), .QN(n4731) );
  NAND3X0 U10079 ( .IN1(n1749), .IN2(g3961), .IN3(g16659), .QN(n4751) );
  NAND3X0 U10080 ( .IN1(g3945), .IN2(n1751), .IN3(g16775), .QN(n4749) );
  NAND3X0 U10081 ( .IN1(n1748), .IN2(g3929), .IN3(g13966), .QN(n4750) );
  NAND3X0 U10082 ( .IN1(n4574), .IN2(n4575), .IN3(n4576), .QN(n4555) );
  NAND3X0 U10083 ( .IN1(n2122), .IN2(g6653), .IN3(g17688), .QN(n4576) );
  NAND3X0 U10084 ( .IN1(g6637), .IN2(n2120), .IN3(g17778), .QN(n4574) );
  NAND3X0 U10085 ( .IN1(n2119), .IN2(g6621), .IN3(g14828), .QN(n4575) );
  NAND3X0 U10086 ( .IN1(n4772), .IN2(n4773), .IN3(n4774), .QN(n4754) );
  NAND3X0 U10087 ( .IN1(n1941), .IN2(g3610), .IN3(g16627), .QN(n4774) );
  NAND3X0 U10088 ( .IN1(g3594), .IN2(n1942), .IN3(g16744), .QN(n4772) );
  NAND3X0 U10089 ( .IN1(n1943), .IN2(g3578), .IN3(g13926), .QN(n4773) );
  NAND3X0 U10090 ( .IN1(n4597), .IN2(n4598), .IN3(n4599), .QN(n4578) );
  NAND3X0 U10091 ( .IN1(n1624), .IN2(g6307), .IN3(g17649), .QN(n4599) );
  NAND3X0 U10092 ( .IN1(g6291), .IN2(n1622), .IN3(g17760), .QN(n4597) );
  NAND3X0 U10093 ( .IN1(n1621), .IN2(g6275), .IN3(g14779), .QN(n4598) );
  NAND3X0 U10094 ( .IN1(g34657), .IN2(n5707), .IN3(g4793), .QN(n4312) );
  NAND3X0 U10095 ( .IN1(g34649), .IN2(n5706), .IN3(g4983), .QN(n4290) );
  NAND3X0 U10096 ( .IN1(n1883), .IN2(g3251), .IN3(g16603), .QN(n4792) );
  NAND3X0 U10097 ( .IN1(n1890), .IN2(g5260), .IN3(g17519), .QN(n4664) );
  NAND3X0 U10098 ( .IN1(n1866), .IN2(g5953), .IN3(g17607), .QN(n4618) );
  NAND3X0 U10099 ( .IN1(n2305), .IN2(g5607), .IN3(g17580), .QN(n4641) );
  NAND3X0 U10100 ( .IN1(n1748), .IN2(g3953), .IN3(g16659), .QN(n4747) );
  NAND3X0 U10101 ( .IN1(n2119), .IN2(g6645), .IN3(g17688), .QN(n4572) );
  NAND3X0 U10102 ( .IN1(n1943), .IN2(test_so43), .IN3(g16627), .QN(n4770) );
  NAND3X0 U10103 ( .IN1(n1621), .IN2(g6299), .IN3(g17649), .QN(n4595) );
  NAND3X0 U10104 ( .IN1(g3235), .IN2(n1880), .IN3(g16718), .QN(n4793) );
  NAND3X0 U10105 ( .IN1(g5244), .IN2(g31860), .IN3(g17674), .QN(n4665) );
  NAND3X0 U10106 ( .IN1(g5937), .IN2(n1870), .IN3(g17739), .QN(n4619) );
  NAND3X0 U10107 ( .IN1(test_so5), .IN2(n2307), .IN3(g17711), .QN(n4642) );
  NAND3X0 U10108 ( .IN1(g3937), .IN2(n1747), .IN3(g16775), .QN(n4748) );
  NAND3X0 U10109 ( .IN1(g6629), .IN2(n2123), .IN3(g17778), .QN(n4573) );
  NAND3X0 U10110 ( .IN1(g3586), .IN2(n1940), .IN3(g16744), .QN(n4771) );
  NAND3X0 U10111 ( .IN1(g6283), .IN2(n1625), .IN3(g17760), .QN(n4596) );
  NAND3X0 U10112 ( .IN1(n2767), .IN2(n2765), .IN3(n4316), .QN(n4315) );
  NAND2X0 U10113 ( .IN1(n2102), .IN2(n5867), .QN(n4316) );
  NBUFFX2 U10114 ( .IN(g1500), .Q(g7946) );
  NBUFFX2 U10115 ( .IN(g1157), .Q(g7916) );
  NAND3X0 U10116 ( .IN1(n4885), .IN2(n5608), .IN3(n4886), .QN(n4882) );
  XNOR2X1 U10117 ( .IN1(g4593), .IN2(g4601), .Q(n4885) );
  XNOR2X1 U10118 ( .IN1(g4584), .IN2(g4608), .Q(n4886) );
  AOI221X1 U10119 ( .IN1(n1880), .IN2(g3347), .IN3(n1881), .IN4(g3343), .IN5(
        n4686), .QN(n4685) );
  OAI22X1 U10120 ( .IN1(g3343), .IN2(n4687), .IN3(g3347), .IN4(n3089), .QN(
        n4686) );
  AOI221X1 U10121 ( .IN1(n1625), .IN2(g6390), .IN3(n1624), .IN4(g6386), .IN5(
        n4696), .QN(n4695) );
  OAI22X1 U10122 ( .IN1(g6386), .IN2(n4589), .IN3(g6390), .IN4(n3028), .QN(
        n4696) );
  AOI221X1 U10123 ( .IN1(n1870), .IN2(test_so50), .IN3(n1869), .IN4(g6040), 
        .IN5(n4702), .QN(n4701) );
  OAI22X1 U10124 ( .IN1(g6040), .IN2(n4612), .IN3(test_so50), .IN4(n3037), 
        .QN(n4702) );
  AOI221X1 U10125 ( .IN1(n1940), .IN2(g3698), .IN3(n1941), .IN4(g3694), .IN5(
        n4681), .QN(n4680) );
  OAI22X1 U10126 ( .IN1(g3694), .IN2(n4682), .IN3(g3698), .IN4(n3078), .QN(
        n4681) );
  AOI221X1 U10127 ( .IN1(n2307), .IN2(g5698), .IN3(n2304), .IN4(g5694), .IN5(
        n4706), .QN(n4705) );
  OAI22X1 U10128 ( .IN1(g5694), .IN2(n4635), .IN3(g5698), .IN4(n3046), .QN(
        n4706) );
  AOI221X1 U10129 ( .IN1(n1747), .IN2(g4049), .IN3(n1749), .IN4(g4045), .IN5(
        n4676), .QN(n4675) );
  OAI22X1 U10130 ( .IN1(g4045), .IN2(n4677), .IN3(g4049), .IN4(n3070), .QN(
        n4676) );
  NOR3X0 U10131 ( .IN1(n5381), .IN2(g1532), .IN3(n5577), .QN(n4894) );
  XOR2X1 U10132 ( .IN1(g239), .IN2(g232), .Q(n5107) );
  OR2X1 U10133 ( .IN1(n2416), .IN2(g2988), .Q(n2778) );
  NAND2X0 U10134 ( .IN1(g1046), .IN2(n1987), .QN(n4807) );
  XNOR2X1 U10135 ( .IN1(n5306), .IN2(g174), .Q(n3679) );
  OA21X1 U10136 ( .IN1(n5265), .IN2(g4366), .IN3(g4369), .Q(g34956) );
  NOR2X0 U10137 ( .IN1(n5266), .IN2(n5267), .QN(n5265) );
  NOR4X0 U10138 ( .IN1(g4311), .IN2(n5540), .IN3(n1492), .IN4(n3094), .QN(
        n5266) );
  NOR4X0 U10139 ( .IN1(n6016), .IN2(g4332), .IN3(g4311), .IN4(n3094), .QN(
        n5267) );
  NOR2X0 U10140 ( .IN1(n6011), .IN2(n6012), .QN(n3282) );
  XOR2X1 U10141 ( .IN1(g4108), .IN2(n6018), .Q(n6011) );
  XOR2X1 U10142 ( .IN1(g4104), .IN2(n6016), .Q(n6012) );
  XNOR2X1 U10143 ( .IN1(g452), .IN2(test_so72), .Q(n3680) );
  OAI22X1 U10144 ( .IN1(n4650), .IN2(n5515), .IN3(g25219), .IN4(n4651), .QN(
        n4649) );
  OA221X1 U10145 ( .IN1(n4652), .IN2(n2739), .IN3(n4653), .IN4(n3056), .IN5(
        n4654), .Q(n4651) );
  OA221X1 U10146 ( .IN1(n4657), .IN2(n4658), .IN3(n5579), .IN4(n4659), .IN5(
        n4660), .Q(n4650) );
  AOI22X1 U10147 ( .IN1(g5208), .IN2(g13039), .IN3(g5220), .IN4(g5339), .QN(
        n4653) );
  AOI22X1 U10148 ( .IN1(g3207), .IN2(g11349), .IN3(g3223), .IN4(g16874), .QN(
        n4781) );
  AOI22X1 U10149 ( .IN1(g5216), .IN2(g12238), .IN3(g5232), .IN4(g17787), .QN(
        n4652) );
  AOI22X1 U10150 ( .IN1(g5909), .IN2(g12350), .IN3(g5925), .IN4(g17819), .QN(
        n4606) );
  AOI22X1 U10151 ( .IN1(g5563), .IN2(g12300), .IN3(g5579), .IN4(g17813), .QN(
        n4629) );
  AOI22X1 U10152 ( .IN1(g3909), .IN2(g11418), .IN3(g3925), .IN4(g16955), .QN(
        n4736) );
  AOI22X1 U10153 ( .IN1(g6601), .IN2(g12470), .IN3(g6617), .IN4(g17871), .QN(
        n4560) );
  AOI22X1 U10154 ( .IN1(g3558), .IN2(g11388), .IN3(g3574), .IN4(g16924), .QN(
        n4759) );
  AOI22X1 U10155 ( .IN1(g6255), .IN2(g12422), .IN3(g6271), .IN4(g17845), .QN(
        n4583) );
  OR2X1 U10156 ( .IN1(n4051), .IN2(test_so53), .Q(n4061) );
  OR2X1 U10157 ( .IN1(n4051), .IN2(g2504), .Q(n4049) );
  NAND2X0 U10158 ( .IN1(n1881), .IN2(g3231), .QN(n4787) );
  NAND2X0 U10159 ( .IN1(n1893), .IN2(g5240), .QN(n4659) );
  NAND2X0 U10160 ( .IN1(n1869), .IN2(g5933), .QN(n4613) );
  NAND2X0 U10161 ( .IN1(n2304), .IN2(g5587), .QN(n4636) );
  NAND2X0 U10162 ( .IN1(n1749), .IN2(g3933), .QN(n4742) );
  NAND2X0 U10163 ( .IN1(n2122), .IN2(g6625), .QN(n4567) );
  NAND2X0 U10164 ( .IN1(n1941), .IN2(g3582), .QN(n4765) );
  NAND2X0 U10165 ( .IN1(n1624), .IN2(g6279), .QN(n4590) );
  NBUFFX2 U10166 ( .IN(g1500), .Q(n6024) );
  NBUFFX2 U10167 ( .IN(g1157), .Q(n6021) );
  AOI22X1 U10168 ( .IN1(g3187), .IN2(g14421), .IN3(test_so88), .IN4(test_so91), 
        .QN(n4786) );
  AOI22X1 U10169 ( .IN1(g5196), .IN2(g13039), .IN3(g5204), .IN4(g5339), .QN(
        n4657) );
  AOI22X1 U10170 ( .IN1(g5889), .IN2(g13068), .IN3(g5897), .IN4(g6031), .QN(
        n4611) );
  AOI22X1 U10171 ( .IN1(g5543), .IN2(g13049), .IN3(g5551), .IN4(g5685), .QN(
        n4634) );
  AOI22X1 U10172 ( .IN1(test_so24), .IN2(g14518), .IN3(g3897), .IN4(g4031), 
        .QN(n4741) );
  AOI22X1 U10173 ( .IN1(g6581), .IN2(g13099), .IN3(g6589), .IN4(g6723), .QN(
        n4565) );
  AOI22X1 U10174 ( .IN1(g3538), .IN2(g14451), .IN3(g3546), .IN4(g3680), .QN(
        n4764) );
  AOI22X1 U10175 ( .IN1(g6235), .IN2(g13085), .IN3(g6243), .IN4(g6377), .QN(
        n4588) );
  OR2X1 U10176 ( .IN1(n5655), .IN2(g1395), .Q(n5217) );
  OR2X1 U10177 ( .IN1(n5654), .IN2(g1052), .Q(n5239) );
  OA22X1 U10178 ( .IN1(n5580), .IN2(n4784), .IN3(n4785), .IN4(n3089), .Q(n4783) );
  NAND2X0 U10179 ( .IN1(n1883), .IN2(g3239), .QN(n4784) );
  AOI22X1 U10180 ( .IN1(g3203), .IN2(g16624), .IN3(g3255), .IN4(g16686), .QN(
        n4785) );
  OA22X1 U10181 ( .IN1(n5579), .IN2(n4655), .IN3(n4656), .IN4(n3055), .Q(n4654) );
  NAND2X0 U10182 ( .IN1(n1890), .IN2(g5248), .QN(n4655) );
  AOI22X1 U10183 ( .IN1(g5212), .IN2(g17577), .IN3(g5264), .IN4(g17639), .QN(
        n4656) );
  OA22X1 U10184 ( .IN1(n5581), .IN2(n4609), .IN3(n4610), .IN4(n3037), .Q(n4608) );
  NAND2X0 U10185 ( .IN1(n1866), .IN2(g5941), .QN(n4609) );
  AOI22X1 U10186 ( .IN1(g5905), .IN2(g17646), .IN3(g5957), .IN4(g17715), .QN(
        n4610) );
  OA22X1 U10187 ( .IN1(n5582), .IN2(n4632), .IN3(n4633), .IN4(n3046), .Q(n4631) );
  NAND2X0 U10188 ( .IN1(n2305), .IN2(g5595), .QN(n4632) );
  AOI22X1 U10189 ( .IN1(test_so6), .IN2(g17604), .IN3(g5611), .IN4(g17678), 
        .QN(n4633) );
  OA22X1 U10190 ( .IN1(n5583), .IN2(n4739), .IN3(n4740), .IN4(n3070), .Q(n4738) );
  NAND2X0 U10191 ( .IN1(n1748), .IN2(g3941), .QN(n4739) );
  AOI22X1 U10192 ( .IN1(g3905), .IN2(g16693), .IN3(g3957), .IN4(g16748), .QN(
        n4740) );
  OA22X1 U10193 ( .IN1(n5584), .IN2(n4563), .IN3(n4564), .IN4(n3017), .Q(n4562) );
  NAND2X0 U10194 ( .IN1(n2119), .IN2(g6633), .QN(n4563) );
  AOI22X1 U10195 ( .IN1(g6597), .IN2(g17722), .IN3(g6649), .IN4(g17764), .QN(
        n4564) );
  OA22X1 U10196 ( .IN1(n5585), .IN2(n4762), .IN3(n4763), .IN4(n3078), .Q(n4761) );
  NAND2X0 U10197 ( .IN1(n1943), .IN2(g3590), .QN(n4762) );
  AOI22X1 U10198 ( .IN1(g3554), .IN2(g16656), .IN3(g3606), .IN4(g16722), .QN(
        n4763) );
  OA22X1 U10199 ( .IN1(n5586), .IN2(n4586), .IN3(n4587), .IN4(n3028), .Q(n4585) );
  NAND2X0 U10200 ( .IN1(n1621), .IN2(g6287), .QN(n4586) );
  AOI22X1 U10201 ( .IN1(g6251), .IN2(g17685), .IN3(g6303), .IN4(g17743), .QN(
        n4587) );
  OAI22X1 U10202 ( .IN1(n4779), .IN2(n5527), .IN3(g3338), .IN4(n4780), .QN(
        n4778) );
  OA221X1 U10203 ( .IN1(n4781), .IN2(n2741), .IN3(n4782), .IN4(n3090), .IN5(
        n4783), .Q(n4780) );
  OA221X1 U10204 ( .IN1(n4786), .IN2(n4687), .IN3(n5580), .IN4(n4787), .IN5(
        n4788), .Q(n4779) );
  AOI22X1 U10205 ( .IN1(g3199), .IN2(g14421), .IN3(g3211), .IN4(test_so91), 
        .QN(n4782) );
  OAI22X1 U10206 ( .IN1(n4604), .IN2(n5528), .IN3(g6035), .IN4(n4605), .QN(
        n4603) );
  OA221X1 U10207 ( .IN1(n4606), .IN2(n2745), .IN3(n4607), .IN4(n3039), .IN5(
        n4608), .Q(n4605) );
  OA221X1 U10208 ( .IN1(n4611), .IN2(n4612), .IN3(n5581), .IN4(n4613), .IN5(
        n4614), .Q(n4604) );
  AOI22X1 U10209 ( .IN1(g5901), .IN2(g13068), .IN3(g5913), .IN4(g6031), .QN(
        n4607) );
  OAI22X1 U10210 ( .IN1(n4627), .IN2(n5529), .IN3(g5689), .IN4(n4628), .QN(
        n4626) );
  OA221X1 U10211 ( .IN1(n4629), .IN2(n2734), .IN3(n4630), .IN4(n3048), .IN5(
        n4631), .Q(n4628) );
  OA221X1 U10212 ( .IN1(n4634), .IN2(n4635), .IN3(n5582), .IN4(n4636), .IN5(
        n4637), .Q(n4627) );
  AOI22X1 U10213 ( .IN1(g5555), .IN2(g13049), .IN3(g5567), .IN4(g5685), .QN(
        n4630) );
  OAI22X1 U10214 ( .IN1(n4734), .IN2(n5530), .IN3(g4040), .IN4(n4735), .QN(
        n4733) );
  OA221X1 U10215 ( .IN1(n4736), .IN2(n2746), .IN3(n4737), .IN4(n3071), .IN5(
        n4738), .Q(n4735) );
  OA221X1 U10216 ( .IN1(n4741), .IN2(n4677), .IN3(n5583), .IN4(n4742), .IN5(
        n4743), .Q(n4734) );
  AOI22X1 U10217 ( .IN1(g3901), .IN2(g14518), .IN3(g3913), .IN4(g4031), .QN(
        n4737) );
  OAI22X1 U10218 ( .IN1(n4558), .IN2(n5531), .IN3(g6727), .IN4(n4559), .QN(
        n4557) );
  OA221X1 U10219 ( .IN1(n4560), .IN2(n2736), .IN3(n4561), .IN4(n3019), .IN5(
        n4562), .Q(n4559) );
  OA221X1 U10220 ( .IN1(n4565), .IN2(n4566), .IN3(n5584), .IN4(n4567), .IN5(
        n4568), .Q(n4558) );
  AOI22X1 U10221 ( .IN1(g6593), .IN2(g13099), .IN3(g6605), .IN4(g6723), .QN(
        n4561) );
  OAI22X1 U10222 ( .IN1(n4757), .IN2(n5532), .IN3(g3689), .IN4(n4758), .QN(
        n4756) );
  OA221X1 U10223 ( .IN1(n4759), .IN2(n2743), .IN3(n4760), .IN4(n3080), .IN5(
        n4761), .Q(n4758) );
  OA221X1 U10224 ( .IN1(n4764), .IN2(n4682), .IN3(n5585), .IN4(n4765), .IN5(
        n4766), .Q(n4757) );
  AOI22X1 U10225 ( .IN1(g3550), .IN2(g14451), .IN3(g3562), .IN4(g3680), .QN(
        n4760) );
  OAI22X1 U10226 ( .IN1(n4581), .IN2(n5533), .IN3(test_so69), .IN4(n4582), 
        .QN(n4580) );
  OA221X1 U10227 ( .IN1(n4583), .IN2(n2742), .IN3(n4584), .IN4(n3029), .IN5(
        n4585), .Q(n4582) );
  OA221X1 U10228 ( .IN1(n4588), .IN2(n4589), .IN3(n5586), .IN4(n4590), .IN5(
        n4591), .Q(n4581) );
  AOI22X1 U10229 ( .IN1(g6247), .IN2(g13085), .IN3(g6259), .IN4(g6377), .QN(
        n4584) );
  NOR4X0 U10230 ( .IN1(n5134), .IN2(g4057), .IN3(g4064), .IN4(g4125), .QN(
        g31521) );
  AND2X1 U10231 ( .IN1(n4724), .IN2(n5135), .Q(n5134) );
  NAND4X0 U10232 ( .IN1(g4112), .IN2(test_so11), .IN3(n1844), .IN4(n5350), 
        .QN(n5135) );
  OAI22X1 U10233 ( .IN1(g6732), .IN2(n4566), .IN3(g6736), .IN4(n3017), .QN(
        n4691) );
  OAI22X1 U10234 ( .IN1(g5348), .IN2(n4658), .IN3(g5352), .IN4(n3055), .QN(
        n4710) );
  NAND4X0 U10235 ( .IN1(n2411), .IN2(n2412), .IN3(n5653), .IN4(n5298), .QN(
        n2410) );
  NAND3X0 U10236 ( .IN1(g4311), .IN2(n5506), .IN3(g4332), .QN(n2412) );
  NAND2X0 U10237 ( .IN1(n2413), .IN2(n5540), .QN(n2411) );
  AO22X1 U10238 ( .IN1(n2414), .IN2(n5506), .IN3(g4322), .IN4(n2415), .Q(n2413) );
  NAND4X0 U10239 ( .IN1(n4287), .IN2(n5713), .IN3(n4288), .IN4(n5318), .QN(
        n4284) );
  NOR2X0 U10240 ( .IN1(g4878), .IN2(g4871), .QN(n4288) );
  NAND4X0 U10241 ( .IN1(n4289), .IN2(n4290), .IN3(n4291), .IN4(n4292), .QN(
        n4287) );
  NAND4X0 U10242 ( .IN1(n4293), .IN2(n5706), .IN3(n5367), .IN4(n5284), .QN(
        n4291) );
  NAND4X0 U10243 ( .IN1(n4309), .IN2(n5712), .IN3(n4310), .IN4(n5440), .QN(
        n4306) );
  NOR2X0 U10244 ( .IN1(g4688), .IN2(g4681), .QN(n4310) );
  NAND4X0 U10245 ( .IN1(n4311), .IN2(n4312), .IN3(n4313), .IN4(n4314), .QN(
        n4309) );
  NAND4X0 U10246 ( .IN1(n4315), .IN2(n5707), .IN3(n5368), .IN4(n5285), .QN(
        n4313) );
  NAND2X0 U10247 ( .IN1(n1864), .IN2(n4058), .QN(n4057) );
  AO221X1 U10248 ( .IN1(n5299), .IN2(n5544), .IN3(g2715), .IN4(n5378), .IN5(
        g2719), .Q(n4058) );
  NAND2X0 U10249 ( .IN1(n1864), .IN2(n4054), .QN(n4053) );
  AO221X1 U10250 ( .IN1(n5299), .IN2(n5545), .IN3(g2715), .IN4(n5379), .IN5(
        g2719), .Q(n4054) );
  INVX0 U10251 ( .IN(g5), .QN(g12833) );
  NAND2X0 U10252 ( .IN1(n4464), .IN2(n4465), .QN(n4463) );
  NAND3X0 U10253 ( .IN1(n5370), .IN2(n5525), .IN3(g1612), .QN(n4465) );
  OR3X1 U10254 ( .IN1(n5587), .IN2(test_so94), .IN3(n5370), .Q(n4464) );
  NAND2X0 U10255 ( .IN1(n4431), .IN2(n4432), .QN(n4430) );
  NAND3X0 U10256 ( .IN1(n5371), .IN2(n5507), .IN3(g2016), .QN(n4432) );
  OR3X1 U10257 ( .IN1(n5683), .IN2(g2051), .IN3(n5371), .Q(n4431) );
  NAND2X0 U10258 ( .IN1(n4453), .IN2(n4454), .QN(n4452) );
  NAND3X0 U10259 ( .IN1(n5602), .IN2(n5359), .IN3(g1748), .QN(n4454) );
  NAND3X0 U10260 ( .IN1(g1752), .IN2(n5596), .IN3(g1760), .QN(n4453) );
  NAND2X0 U10261 ( .IN1(n4385), .IN2(n4386), .QN(n4384) );
  NAND3X0 U10262 ( .IN1(n5372), .IN2(n5508), .IN3(test_so66), .QN(n4386) );
  OR3X1 U10263 ( .IN1(n5684), .IN2(g2610), .IN3(n5372), .Q(n4385) );
  NAND2X0 U10264 ( .IN1(n4397), .IN2(n4398), .QN(n4396) );
  NAND3X0 U10265 ( .IN1(n5373), .IN2(n5509), .IN3(g2441), .QN(n4398) );
  OR3X1 U10266 ( .IN1(n5685), .IN2(g2476), .IN3(n5373), .Q(n4397) );
  NAND2X0 U10267 ( .IN1(n4442), .IN2(n4443), .QN(n4441) );
  NAND3X0 U10268 ( .IN1(n5374), .IN2(n5510), .IN3(g1882), .QN(n4443) );
  OR3X1 U10269 ( .IN1(n5686), .IN2(g1917), .IN3(n5374), .Q(n4442) );
  NAND2X0 U10270 ( .IN1(n4408), .IN2(n4409), .QN(n4407) );
  NAND3X0 U10271 ( .IN1(n5375), .IN2(n5511), .IN3(g2307), .QN(n4409) );
  OR3X1 U10272 ( .IN1(n5687), .IN2(test_so21), .IN3(n5375), .Q(n4408) );
  NAND2X0 U10273 ( .IN1(n4420), .IN2(n4421), .QN(n4419) );
  NAND3X0 U10274 ( .IN1(n5376), .IN2(n5512), .IN3(g2173), .QN(n4421) );
  OR3X1 U10275 ( .IN1(n5688), .IN2(g2208), .IN3(n5376), .Q(n4420) );
  NAND2X0 U10276 ( .IN1(g4515), .IN2(n1490), .QN(n2415) );
  NAND3X0 U10277 ( .IN1(n2752), .IN2(n2750), .IN3(n4294), .QN(n4293) );
  NAND2X0 U10278 ( .IN1(n2134), .IN2(n5879), .QN(n4294) );
  NAND2X0 U10279 ( .IN1(g1442), .IN2(n5617), .QN(n4899) );
  NAND2X0 U10280 ( .IN1(g3863), .IN2(g3857), .QN(n3479) );
  NAND2X0 U10281 ( .IN1(g6555), .IN2(g6549), .QN(n3404) );
  NAND2X0 U10282 ( .IN1(g5863), .IN2(g5857), .QN(n3424) );
  NAND2X0 U10283 ( .IN1(g5170), .IN2(g5164), .QN(n3444) );
  NAND2X0 U10284 ( .IN1(g6209), .IN2(g6203), .QN(n3414) );
  NAND2X0 U10285 ( .IN1(g3512), .IN2(g3506), .QN(n3489) );
  NAND2X0 U10286 ( .IN1(g5517), .IN2(g5511), .QN(n3434) );
  NAND2X0 U10287 ( .IN1(g3161), .IN2(g3155), .QN(n3500) );
  NAND2X0 U10288 ( .IN1(test_so7), .IN2(n5618), .QN(n4924) );
  NAND2X0 U10289 ( .IN1(n1732), .IN2(g3167), .QN(n3496) );
  OA22X1 U10290 ( .IN1(n5317), .IN2(g324), .IN3(n5827), .IN4(n5282), .Q(n4971)
         );
  NOR2X0 U10291 ( .IN1(g355), .IN2(g333), .QN(n4966) );
  NOR2X0 U10292 ( .IN1(test_so7), .IN2(g1146), .QN(n4496) );
  NOR2X0 U10293 ( .IN1(g1442), .IN2(g1489), .QN(n4472) );
  NAND2X0 U10294 ( .IN1(g218), .IN2(g8291), .QN(n5131) );
  AND4X1 U10295 ( .IN1(DFF_348_n1), .IN2(n5819), .IN3(DFF_1225_n1), .IN4(n4867), .Q(n4861) );
  NOR2X0 U10296 ( .IN1(test_so47), .IN2(g4438), .QN(n4867) );
  NAND2X0 U10297 ( .IN1(g5170), .IN2(n5570), .QN(n3446) );
  NAND2X0 U10298 ( .IN1(g6555), .IN2(n5571), .QN(n3406) );
  NAND2X0 U10299 ( .IN1(g3863), .IN2(n5572), .QN(n3481) );
  NAND2X0 U10300 ( .IN1(g5863), .IN2(n5573), .QN(n3426) );
  NAND2X0 U10301 ( .IN1(g6209), .IN2(n5574), .QN(n3416) );
  NAND2X0 U10302 ( .IN1(g5517), .IN2(n5575), .QN(n3436) );
  NAND2X0 U10303 ( .IN1(g3512), .IN2(n5576), .QN(n3491) );
  NAND2X0 U10304 ( .IN1(g3161), .IN2(n5366), .QN(n3502) );
  NAND2X0 U10305 ( .IN1(g1105), .IN2(n4492), .QN(n4931) );
  AND4X1 U10306 ( .IN1(g4492), .IN2(g4489), .IN3(test_so27), .IN4(g4483), .Q(
        n2777) );
  NAND2X0 U10307 ( .IN1(g1448), .IN2(n4468), .QN(n4906) );
  NAND3X0 U10308 ( .IN1(test_so3), .IN2(n5727), .IN3(g4633), .QN(n4880) );
  NAND2X0 U10309 ( .IN1(g812), .IN2(g847), .QN(n5244) );
  NAND2X0 U10310 ( .IN1(g817), .IN2(n5709), .QN(n5247) );
  OR2X1 U10311 ( .IN1(n5366), .IN2(g3161), .Q(n3501) );
  NAND2X0 U10312 ( .IN1(n2563), .IN2(g4849), .QN(n2561) );
  NAND2X0 U10313 ( .IN1(n2573), .IN2(g4659), .QN(n2571) );
  ISOLANDX1 U10314 ( .D(g667), .ISO(g686), .Q(n4962) );
  NAND2X0 U10315 ( .IN1(g827), .IN2(g832), .QN(n5243) );
  NAND3X0 U10316 ( .IN1(g1548), .IN2(g1430), .IN3(g1564), .QN(n5049) );
  NAND3X0 U10317 ( .IN1(g1205), .IN2(g1087), .IN3(g1221), .QN(n5075) );
  ISOLANDX1 U10318 ( .D(g5092), .ISO(n5681), .Q(n5016) );
  NAND3X0 U10319 ( .IN1(n5682), .IN2(n5431), .IN3(g890), .QN(n4946) );
  XOR2X1 U10320 ( .IN1(g9251), .IN2(g4308), .Q(n5168) );
  XOR2X1 U10321 ( .IN1(g9019), .IN2(g4291), .Q(n5258) );
  XOR2X1 U10322 ( .IN1(g8839), .IN2(g4281), .Q(n5260) );
  XOR2X1 U10323 ( .IN1(n2777), .IN2(g4527), .Q(n4713) );
  OAI22X1 U10324 ( .IN1(n5484), .IN2(g4164), .IN3(g4145), .IN4(g4253), .QN(
        n5175) );

  HighActiveRegionDetection TrojanTrigger (CK, g26963, g34629, g25757, g34640, g34628, g26888, g34635, g34619, Tj_Trigger); 
  
  // When the Trojan is triggered, it leaks the value of g25715 signal through g10122_Tj output pin.
   MUX21X1 Trojan_Paylod ( .IN1(g10122_Tj), .IN2(g25715), .S(Trigger_out), .Q(g10122) );
endmodule

